magic
tech sky130A
timestamp 1634770709
<< nmos >>
rect 340 155 840 205
rect 340 55 840 105
<< ndiff >>
rect 340 240 840 250
rect 340 220 355 240
rect 375 220 395 240
rect 415 220 435 240
rect 455 220 475 240
rect 495 220 515 240
rect 535 220 555 240
rect 575 220 595 240
rect 615 220 635 240
rect 655 220 675 240
rect 695 220 715 240
rect 735 220 755 240
rect 775 220 795 240
rect 825 220 840 240
rect 340 205 840 220
rect 340 140 840 155
rect 340 120 355 140
rect 375 120 395 140
rect 415 120 435 140
rect 455 120 475 140
rect 495 120 515 140
rect 535 120 555 140
rect 575 120 595 140
rect 615 120 635 140
rect 655 120 675 140
rect 695 120 715 140
rect 735 120 755 140
rect 775 120 795 140
rect 825 120 840 140
rect 340 105 840 120
rect 340 40 840 55
rect 340 20 355 40
rect 375 20 395 40
rect 415 20 435 40
rect 455 20 475 40
rect 495 20 515 40
rect 535 20 555 40
rect 575 20 595 40
rect 615 20 635 40
rect 655 20 675 40
rect 695 20 715 40
rect 735 20 755 40
rect 775 20 795 40
rect 825 20 840 40
rect 340 10 840 20
<< ndiffc >>
rect 355 220 375 240
rect 395 220 415 240
rect 435 220 455 240
rect 475 220 495 240
rect 515 220 535 240
rect 555 220 575 240
rect 595 220 615 240
rect 635 220 655 240
rect 675 220 695 240
rect 715 220 735 240
rect 755 220 775 240
rect 795 220 825 240
rect 355 120 375 140
rect 395 120 415 140
rect 435 120 455 140
rect 475 120 495 140
rect 515 120 535 140
rect 555 120 575 140
rect 595 120 615 140
rect 635 120 655 140
rect 675 120 695 140
rect 715 120 735 140
rect 755 120 775 140
rect 795 120 825 140
rect 355 20 375 40
rect 395 20 415 40
rect 435 20 455 40
rect 475 20 495 40
rect 515 20 535 40
rect 555 20 575 40
rect 595 20 615 40
rect 635 20 655 40
rect 675 20 695 40
rect 715 20 735 40
rect 755 20 775 40
rect 795 20 825 40
<< psubdiff >>
rect 340 280 840 290
rect 340 260 355 280
rect 375 260 395 280
rect 415 260 435 280
rect 455 260 475 280
rect 495 260 515 280
rect 535 260 555 280
rect 575 260 595 280
rect 615 260 635 280
rect 655 260 675 280
rect 695 260 715 280
rect 735 260 755 280
rect 775 260 795 280
rect 825 260 840 280
rect 340 250 840 260
<< psubdiffcont >>
rect 355 260 375 280
rect 395 260 415 280
rect 435 260 455 280
rect 475 260 495 280
rect 515 260 535 280
rect 555 260 575 280
rect 595 260 615 280
rect 635 260 655 280
rect 675 260 695 280
rect 715 260 735 280
rect 755 260 775 280
rect 795 260 825 280
<< poly >>
rect 325 155 340 205
rect 840 195 900 205
rect 840 165 870 195
rect 890 165 900 195
rect 840 155 900 165
rect 325 55 340 105
rect 840 95 900 105
rect 840 65 870 95
rect 890 65 900 95
rect 840 55 900 65
<< polycont >>
rect 870 165 890 195
rect 870 65 890 95
<< xpolycontact >>
rect 950 1610 1170 1645
rect 2770 1610 2990 1645
rect 950 1450 1170 1485
rect 2770 1450 2990 1485
rect 950 1290 1170 1325
rect 2770 1290 2990 1325
rect 950 1130 1170 1165
rect 2770 1130 2990 1165
rect 950 970 1170 1005
rect 2770 970 2990 1005
rect 950 810 1170 845
rect 2770 810 2990 845
rect 950 650 1170 685
rect 2770 650 2990 685
rect 950 490 1170 525
rect 2770 490 2990 525
rect 950 330 1170 365
rect 2770 330 2990 365
rect 950 170 1170 205
rect 2770 170 2990 205
rect 950 10 1170 45
rect 2770 10 2990 45
<< xpolyres >>
rect 1170 1610 2770 1645
rect 1170 1450 2770 1485
rect 1170 1290 2770 1325
rect 1170 1130 2770 1165
rect 1170 970 2770 1005
rect 1170 810 2770 845
rect 1170 650 2770 685
rect 1170 490 2770 525
rect 1170 330 2770 365
rect 1170 170 2770 205
rect 1170 10 2770 45
<< locali >>
rect 340 280 840 290
rect 340 260 355 280
rect 375 260 395 280
rect 415 260 435 280
rect 455 260 475 280
rect 495 260 515 280
rect 535 260 555 280
rect 575 260 595 280
rect 615 260 635 280
rect 655 260 675 280
rect 695 260 715 280
rect 735 260 755 280
rect 775 260 795 280
rect 825 260 840 280
rect 340 240 840 260
rect 340 220 355 240
rect 375 220 395 240
rect 415 220 435 240
rect 455 220 475 240
rect 495 220 515 240
rect 535 220 555 240
rect 575 220 595 240
rect 615 220 635 240
rect 655 220 675 240
rect 695 220 715 240
rect 735 220 755 240
rect 775 220 795 240
rect 825 220 840 240
rect 340 210 840 220
rect 860 195 900 205
rect 860 165 870 195
rect 890 165 900 195
rect 860 150 900 165
rect 340 145 900 150
rect 340 140 870 145
rect 340 120 355 140
rect 375 120 395 140
rect 415 120 435 140
rect 455 120 475 140
rect 495 120 515 140
rect 535 120 555 140
rect 575 120 595 140
rect 615 120 635 140
rect 655 120 675 140
rect 695 120 715 140
rect 735 120 755 140
rect 775 120 795 140
rect 825 120 870 140
rect 340 115 870 120
rect 890 115 900 145
rect 340 110 900 115
rect 860 95 900 110
rect 860 65 870 95
rect 890 65 900 95
rect 860 55 900 65
rect 340 40 840 50
rect 340 20 355 40
rect 375 20 395 40
rect 415 20 435 40
rect 455 20 475 40
rect 495 20 515 40
rect 535 20 555 40
rect 575 20 595 40
rect 615 20 635 40
rect 655 20 675 40
rect 695 20 715 40
rect 735 20 755 40
rect 775 20 795 40
rect 825 20 840 40
rect 340 10 840 20
<< viali >>
rect 980 1615 1000 1640
rect 1020 1615 1040 1640
rect 1060 1615 1080 1640
rect 1100 1615 1120 1640
rect 1140 1615 1160 1640
rect 2780 1615 2800 1640
rect 2820 1615 2840 1640
rect 2860 1615 2880 1640
rect 2900 1615 2920 1640
rect 2940 1615 2960 1640
rect 980 1455 1000 1480
rect 1020 1455 1040 1480
rect 1060 1455 1080 1480
rect 1100 1455 1120 1480
rect 1140 1455 1160 1480
rect 2780 1455 2800 1480
rect 2820 1455 2840 1480
rect 2860 1455 2880 1480
rect 2900 1455 2920 1480
rect 2940 1455 2960 1480
rect 980 1295 1000 1320
rect 1020 1295 1040 1320
rect 1060 1295 1080 1320
rect 1100 1295 1120 1320
rect 1140 1295 1160 1320
rect 2780 1295 2800 1320
rect 2820 1295 2840 1320
rect 2860 1295 2880 1320
rect 2900 1295 2920 1320
rect 2940 1295 2960 1320
rect 980 1135 1000 1160
rect 1020 1135 1040 1160
rect 1060 1135 1080 1160
rect 1100 1135 1120 1160
rect 1140 1135 1160 1160
rect 2780 1135 2800 1160
rect 2820 1135 2840 1160
rect 2860 1135 2880 1160
rect 2900 1135 2920 1160
rect 2940 1135 2960 1160
rect 980 975 1000 1000
rect 1020 975 1040 1000
rect 1060 975 1080 1000
rect 1100 975 1120 1000
rect 1140 975 1160 1000
rect 2780 975 2800 1000
rect 2820 975 2840 1000
rect 2860 975 2880 1000
rect 2900 975 2920 1000
rect 2940 975 2960 1000
rect 980 815 1000 840
rect 1020 815 1040 840
rect 1060 815 1080 840
rect 1100 815 1120 840
rect 1140 815 1160 840
rect 2780 815 2800 840
rect 2820 815 2840 840
rect 2860 815 2880 840
rect 2900 815 2920 840
rect 2940 815 2960 840
rect 980 655 1000 680
rect 1020 655 1040 680
rect 1060 655 1080 680
rect 1100 655 1120 680
rect 1140 655 1160 680
rect 2780 655 2800 680
rect 2820 655 2840 680
rect 2860 655 2880 680
rect 2900 655 2920 680
rect 2940 655 2960 680
rect 980 495 1000 520
rect 1020 495 1040 520
rect 1060 495 1080 520
rect 1100 495 1120 520
rect 1140 495 1160 520
rect 2780 495 2800 520
rect 2820 495 2840 520
rect 2860 495 2880 520
rect 2900 495 2920 520
rect 2940 495 2960 520
rect 980 335 1000 360
rect 1020 335 1040 360
rect 1060 335 1080 360
rect 1100 335 1120 360
rect 1140 335 1160 360
rect 2780 335 2800 360
rect 2820 335 2840 360
rect 2860 335 2880 360
rect 2900 335 2920 360
rect 2940 335 2960 360
rect 355 260 375 280
rect 395 260 415 280
rect 435 260 455 280
rect 475 260 495 280
rect 515 260 535 280
rect 555 260 575 280
rect 595 260 615 280
rect 635 260 655 280
rect 675 260 695 280
rect 715 260 735 280
rect 755 260 775 280
rect 795 260 825 280
rect 355 220 375 240
rect 395 220 415 240
rect 435 220 455 240
rect 475 220 495 240
rect 515 220 535 240
rect 555 220 575 240
rect 595 220 615 240
rect 635 220 655 240
rect 675 220 695 240
rect 715 220 735 240
rect 755 220 775 240
rect 795 220 825 240
rect 870 165 890 195
rect 980 175 1000 200
rect 1020 175 1040 200
rect 1060 175 1080 200
rect 1100 175 1120 200
rect 1140 175 1160 200
rect 2780 175 2800 200
rect 2820 175 2840 200
rect 2860 175 2880 200
rect 2900 175 2920 200
rect 2940 175 2960 200
rect 355 120 375 140
rect 395 120 415 140
rect 435 120 455 140
rect 475 120 495 140
rect 515 120 535 140
rect 555 120 575 140
rect 595 120 615 140
rect 635 120 655 140
rect 675 120 695 140
rect 715 120 735 140
rect 755 120 775 140
rect 795 120 825 140
rect 870 115 890 145
rect 870 65 890 95
rect 355 20 375 40
rect 395 20 415 40
rect 435 20 455 40
rect 475 20 495 40
rect 515 20 535 40
rect 555 20 575 40
rect 595 20 615 40
rect 635 20 655 40
rect 675 20 695 40
rect 715 20 735 40
rect 755 20 775 40
rect 795 20 825 40
rect 980 15 1000 40
rect 1020 15 1040 40
rect 1060 15 1080 40
rect 1100 15 1120 40
rect 1140 15 1160 40
rect 2780 15 2800 40
rect 2820 15 2840 40
rect 2860 15 2880 40
rect 2900 15 2920 40
rect 2940 15 2960 40
<< metal1 >>
rect 950 1640 1170 1645
rect 950 1615 980 1640
rect 1000 1615 1020 1640
rect 1040 1615 1060 1640
rect 1080 1615 1100 1640
rect 1120 1615 1140 1640
rect 1160 1615 1170 1640
rect 950 1480 1170 1615
rect 2770 1640 2990 1645
rect 2770 1610 2780 1640
rect 2810 1610 2820 1640
rect 2850 1610 2860 1640
rect 2890 1610 2900 1640
rect 2930 1610 2940 1640
rect 2970 1610 2990 1640
rect 950 1455 980 1480
rect 1000 1455 1020 1480
rect 1040 1455 1060 1480
rect 1080 1455 1100 1480
rect 1120 1455 1140 1480
rect 1160 1455 1170 1480
rect 950 1450 1170 1455
rect 2770 1480 2990 1485
rect 2770 1455 2780 1480
rect 2800 1455 2820 1480
rect 2840 1455 2860 1480
rect 2880 1455 2900 1480
rect 2920 1455 2940 1480
rect 2960 1455 2990 1480
rect 950 1320 1170 1325
rect 950 1295 980 1320
rect 1000 1295 1020 1320
rect 1040 1295 1060 1320
rect 1080 1295 1100 1320
rect 1120 1295 1140 1320
rect 1160 1295 1170 1320
rect 950 1160 1170 1295
rect 2770 1320 2990 1455
rect 2770 1295 2780 1320
rect 2800 1295 2820 1320
rect 2840 1295 2860 1320
rect 2880 1295 2900 1320
rect 2920 1295 2940 1320
rect 2960 1295 2990 1320
rect 2770 1290 2990 1295
rect 950 1135 980 1160
rect 1000 1135 1020 1160
rect 1040 1135 1060 1160
rect 1080 1135 1100 1160
rect 1120 1135 1140 1160
rect 1160 1135 1170 1160
rect 950 1130 1170 1135
rect 2770 1160 2990 1165
rect 2770 1135 2780 1160
rect 2800 1135 2820 1160
rect 2840 1135 2860 1160
rect 2880 1135 2900 1160
rect 2920 1135 2940 1160
rect 2960 1135 2990 1160
rect 950 1000 1170 1005
rect 950 975 980 1000
rect 1000 975 1020 1000
rect 1040 975 1060 1000
rect 1080 975 1100 1000
rect 1120 975 1140 1000
rect 1160 975 1170 1000
rect 950 840 1170 975
rect 2770 1000 2990 1135
rect 2770 975 2780 1000
rect 2800 975 2820 1000
rect 2840 975 2860 1000
rect 2880 975 2900 1000
rect 2920 975 2940 1000
rect 2960 975 2990 1000
rect 2770 970 2990 975
rect 950 815 980 840
rect 1000 815 1020 840
rect 1040 815 1060 840
rect 1080 815 1100 840
rect 1120 815 1140 840
rect 1160 815 1170 840
rect 950 810 1170 815
rect 2770 840 2990 845
rect 2770 815 2780 840
rect 2800 815 2820 840
rect 2840 815 2860 840
rect 2880 815 2900 840
rect 2920 815 2940 840
rect 2960 815 2990 840
rect 950 680 1170 685
rect 950 655 980 680
rect 1000 655 1020 680
rect 1040 655 1060 680
rect 1080 655 1100 680
rect 1120 655 1140 680
rect 1160 655 1170 680
rect 950 520 1170 655
rect 2770 680 2990 815
rect 2770 655 2780 680
rect 2800 655 2820 680
rect 2840 655 2860 680
rect 2880 655 2900 680
rect 2920 655 2940 680
rect 2960 655 2990 680
rect 2770 650 2990 655
rect 950 495 980 520
rect 1000 495 1020 520
rect 1040 495 1060 520
rect 1080 495 1100 520
rect 1120 495 1140 520
rect 1160 495 1170 520
rect 950 490 1170 495
rect 2770 520 2990 525
rect 2770 495 2780 520
rect 2800 495 2820 520
rect 2840 495 2860 520
rect 2880 495 2900 520
rect 2920 495 2940 520
rect 2960 495 2990 520
rect 950 360 1170 365
rect 950 335 980 360
rect 1000 335 1020 360
rect 1040 335 1060 360
rect 1080 335 1100 360
rect 1120 335 1140 360
rect 1160 335 1170 360
rect 340 280 840 290
rect 340 260 355 280
rect 375 260 395 280
rect 415 260 435 280
rect 455 260 475 280
rect 495 260 515 280
rect 535 260 555 280
rect 575 260 595 280
rect 615 260 635 280
rect 655 260 675 280
rect 695 260 715 280
rect 735 260 755 280
rect 775 260 795 280
rect 825 260 840 280
rect 340 240 840 260
rect 340 220 355 240
rect 375 220 395 240
rect 415 220 435 240
rect 455 220 475 240
rect 495 220 515 240
rect 535 220 555 240
rect 575 220 595 240
rect 615 220 635 240
rect 655 220 675 240
rect 695 220 715 240
rect 735 220 755 240
rect 775 220 795 240
rect 825 220 840 240
rect 340 210 840 220
rect 860 195 900 205
rect 860 165 870 195
rect 890 165 900 195
rect 950 200 1170 335
rect 2770 360 2990 495
rect 2770 335 2780 360
rect 2800 335 2820 360
rect 2840 335 2860 360
rect 2880 335 2900 360
rect 2920 335 2940 360
rect 2960 335 2990 360
rect 2770 330 2990 335
rect 950 175 980 200
rect 1000 175 1020 200
rect 1040 175 1060 200
rect 1080 175 1100 200
rect 1120 175 1140 200
rect 1160 175 1170 200
rect 950 170 1170 175
rect 2770 200 2990 205
rect 2770 175 2780 200
rect 2800 175 2820 200
rect 2840 175 2860 200
rect 2880 175 2900 200
rect 2920 175 2940 200
rect 2960 175 2990 200
rect 340 140 840 150
rect 340 120 355 140
rect 375 120 395 140
rect 415 120 435 140
rect 455 120 475 140
rect 495 120 515 140
rect 535 120 555 140
rect 575 120 595 140
rect 615 120 635 140
rect 655 120 675 140
rect 695 120 715 140
rect 735 120 755 140
rect 775 120 795 140
rect 825 120 840 140
rect 340 110 840 120
rect 860 145 900 165
rect 860 115 870 145
rect 890 115 900 145
rect 860 95 900 115
rect 860 65 870 95
rect 890 65 900 95
rect 340 40 840 50
rect 340 20 355 40
rect 375 20 395 40
rect 415 20 435 40
rect 455 20 475 40
rect 495 20 515 40
rect 535 20 555 40
rect 575 20 595 40
rect 615 20 635 40
rect 655 20 675 40
rect 695 20 715 40
rect 735 20 755 40
rect 775 20 795 40
rect 825 20 840 40
rect 340 10 840 20
rect 860 45 900 65
rect 860 40 1170 45
rect 860 15 980 40
rect 1000 15 1020 40
rect 1040 15 1060 40
rect 1080 15 1100 40
rect 1120 15 1140 40
rect 1160 15 1170 40
rect 860 10 1170 15
rect 2770 40 2990 175
rect 2770 15 2780 40
rect 2800 15 2820 40
rect 2840 15 2860 40
rect 2880 15 2900 40
rect 2920 15 2940 40
rect 2960 15 2990 40
rect 2770 10 2990 15
<< via1 >>
rect 2780 1615 2800 1640
rect 2800 1615 2810 1640
rect 2780 1610 2810 1615
rect 2820 1615 2840 1640
rect 2840 1615 2850 1640
rect 2820 1610 2850 1615
rect 2860 1615 2880 1640
rect 2880 1615 2890 1640
rect 2860 1610 2890 1615
rect 2900 1615 2920 1640
rect 2920 1615 2930 1640
rect 2900 1610 2930 1615
rect 2940 1615 2960 1640
rect 2960 1615 2970 1640
rect 2940 1610 2970 1615
<< metal2 >>
rect 2770 1640 2990 1645
rect 2770 1610 2780 1640
rect 2810 1610 2820 1640
rect 2855 1610 2860 1640
rect 2970 1610 2990 1640
rect 2770 1605 2990 1610
<< via2 >>
rect 2780 1610 2810 1640
rect 2825 1610 2850 1640
rect 2850 1610 2855 1640
rect 2870 1610 2890 1640
rect 2890 1610 2900 1640
rect 2915 1610 2930 1640
rect 2930 1610 2940 1640
rect 2940 1610 2945 1640
<< metal3 >>
rect 2770 1640 2970 1645
rect 2770 1605 2780 1640
rect 2815 1610 2825 1640
rect 2865 1610 2870 1640
rect 2815 1605 2830 1610
rect 2865 1605 2880 1610
rect 2915 1605 2930 1610
rect 2965 1605 2970 1640
rect 3010 -130 4620 1645
rect 3010 -165 3030 -130
rect 3065 -165 3075 -130
rect 3110 -165 3120 -130
rect 3155 -165 3165 -130
rect 3200 -165 3210 -130
rect 3245 -165 3255 -130
rect 3290 -165 3300 -130
rect 3335 -165 3345 -130
rect 3380 -165 3390 -130
rect 3425 -165 3435 -130
rect 3470 -165 3480 -130
rect 3515 -165 3525 -130
rect 3560 -165 3570 -130
rect 3605 -165 3615 -130
rect 3650 -165 3660 -130
rect 3695 -165 3705 -130
rect 3740 -165 3750 -130
rect 3785 -165 3795 -130
rect 3830 -165 3840 -130
rect 3875 -165 3885 -130
rect 3920 -165 3930 -130
rect 3965 -165 3975 -130
rect 4010 -165 4020 -130
rect 4055 -165 4065 -130
rect 4100 -165 4110 -130
rect 4145 -165 4155 -130
rect 4190 -165 4200 -130
rect 4235 -165 4245 -130
rect 4280 -165 4290 -130
rect 4325 -165 4335 -130
rect 4370 -165 4380 -130
rect 4415 -165 4425 -130
rect 4460 -165 4470 -130
rect 4505 -165 4515 -130
rect 4550 -165 4560 -130
rect 4595 -165 4620 -130
rect 3010 -175 4620 -165
rect 3010 -210 3030 -175
rect 3065 -210 3075 -175
rect 3110 -210 3120 -175
rect 3155 -210 3165 -175
rect 3200 -210 3210 -175
rect 3245 -210 3255 -175
rect 3290 -210 3300 -175
rect 3335 -210 3345 -175
rect 3380 -210 3390 -175
rect 3425 -210 3435 -175
rect 3470 -210 3480 -175
rect 3515 -210 3525 -175
rect 3560 -210 3570 -175
rect 3605 -210 3615 -175
rect 3650 -210 3660 -175
rect 3695 -210 3705 -175
rect 3740 -210 3750 -175
rect 3785 -210 3795 -175
rect 3830 -210 3840 -175
rect 3875 -210 3885 -175
rect 3920 -210 3930 -175
rect 3965 -210 3975 -175
rect 4010 -210 4020 -175
rect 4055 -210 4065 -175
rect 4100 -210 4110 -175
rect 4145 -210 4155 -175
rect 4190 -210 4200 -175
rect 4235 -210 4245 -175
rect 4280 -210 4290 -175
rect 4325 -210 4335 -175
rect 4370 -210 4380 -175
rect 4415 -210 4425 -175
rect 4460 -210 4470 -175
rect 4505 -210 4515 -175
rect 4550 -210 4560 -175
rect 4595 -210 4620 -175
rect 3010 -220 4620 -210
rect 3010 -255 3030 -220
rect 3065 -255 3075 -220
rect 3110 -255 3120 -220
rect 3155 -255 3165 -220
rect 3200 -255 3210 -220
rect 3245 -255 3255 -220
rect 3290 -255 3300 -220
rect 3335 -255 3345 -220
rect 3380 -255 3390 -220
rect 3425 -255 3435 -220
rect 3470 -255 3480 -220
rect 3515 -255 3525 -220
rect 3560 -255 3570 -220
rect 3605 -255 3615 -220
rect 3650 -255 3660 -220
rect 3695 -255 3705 -220
rect 3740 -255 3750 -220
rect 3785 -255 3795 -220
rect 3830 -255 3840 -220
rect 3875 -255 3885 -220
rect 3920 -255 3930 -220
rect 3965 -255 3975 -220
rect 4010 -255 4020 -220
rect 4055 -255 4065 -220
rect 4100 -255 4110 -220
rect 4145 -255 4155 -220
rect 4190 -255 4200 -220
rect 4235 -255 4245 -220
rect 4280 -255 4290 -220
rect 4325 -255 4335 -220
rect 4370 -255 4380 -220
rect 4415 -255 4425 -220
rect 4460 -255 4470 -220
rect 4505 -255 4515 -220
rect 4550 -255 4560 -220
rect 4595 -255 4620 -220
rect 3010 -285 4620 -255
<< via3 >>
rect 2780 1610 2810 1640
rect 2810 1610 2815 1640
rect 2830 1610 2855 1640
rect 2855 1610 2865 1640
rect 2880 1610 2900 1640
rect 2900 1610 2915 1640
rect 2930 1610 2945 1640
rect 2945 1610 2965 1640
rect 2780 1605 2815 1610
rect 2830 1605 2865 1610
rect 2880 1605 2915 1610
rect 2930 1605 2965 1610
rect 3030 -165 3065 -130
rect 3075 -165 3110 -130
rect 3120 -165 3155 -130
rect 3165 -165 3200 -130
rect 3210 -165 3245 -130
rect 3255 -165 3290 -130
rect 3300 -165 3335 -130
rect 3345 -165 3380 -130
rect 3390 -165 3425 -130
rect 3435 -165 3470 -130
rect 3480 -165 3515 -130
rect 3525 -165 3560 -130
rect 3570 -165 3605 -130
rect 3615 -165 3650 -130
rect 3660 -165 3695 -130
rect 3705 -165 3740 -130
rect 3750 -165 3785 -130
rect 3795 -165 3830 -130
rect 3840 -165 3875 -130
rect 3885 -165 3920 -130
rect 3930 -165 3965 -130
rect 3975 -165 4010 -130
rect 4020 -165 4055 -130
rect 4065 -165 4100 -130
rect 4110 -165 4145 -130
rect 4155 -165 4190 -130
rect 4200 -165 4235 -130
rect 4245 -165 4280 -130
rect 4290 -165 4325 -130
rect 4335 -165 4370 -130
rect 4380 -165 4415 -130
rect 4425 -165 4460 -130
rect 4470 -165 4505 -130
rect 4515 -165 4550 -130
rect 4560 -165 4595 -130
rect 3030 -210 3065 -175
rect 3075 -210 3110 -175
rect 3120 -210 3155 -175
rect 3165 -210 3200 -175
rect 3210 -210 3245 -175
rect 3255 -210 3290 -175
rect 3300 -210 3335 -175
rect 3345 -210 3380 -175
rect 3390 -210 3425 -175
rect 3435 -210 3470 -175
rect 3480 -210 3515 -175
rect 3525 -210 3560 -175
rect 3570 -210 3605 -175
rect 3615 -210 3650 -175
rect 3660 -210 3695 -175
rect 3705 -210 3740 -175
rect 3750 -210 3785 -175
rect 3795 -210 3830 -175
rect 3840 -210 3875 -175
rect 3885 -210 3920 -175
rect 3930 -210 3965 -175
rect 3975 -210 4010 -175
rect 4020 -210 4055 -175
rect 4065 -210 4100 -175
rect 4110 -210 4145 -175
rect 4155 -210 4190 -175
rect 4200 -210 4235 -175
rect 4245 -210 4280 -175
rect 4290 -210 4325 -175
rect 4335 -210 4370 -175
rect 4380 -210 4415 -175
rect 4425 -210 4460 -175
rect 4470 -210 4505 -175
rect 4515 -210 4550 -175
rect 4560 -210 4595 -175
rect 3030 -255 3065 -220
rect 3075 -255 3110 -220
rect 3120 -255 3155 -220
rect 3165 -255 3200 -220
rect 3210 -255 3245 -220
rect 3255 -255 3290 -220
rect 3300 -255 3335 -220
rect 3345 -255 3380 -220
rect 3390 -255 3425 -220
rect 3435 -255 3470 -220
rect 3480 -255 3515 -220
rect 3525 -255 3560 -220
rect 3570 -255 3605 -220
rect 3615 -255 3650 -220
rect 3660 -255 3695 -220
rect 3705 -255 3740 -220
rect 3750 -255 3785 -220
rect 3795 -255 3830 -220
rect 3840 -255 3875 -220
rect 3885 -255 3920 -220
rect 3930 -255 3965 -220
rect 3975 -255 4010 -220
rect 4020 -255 4055 -220
rect 4065 -255 4100 -220
rect 4110 -255 4145 -220
rect 4155 -255 4190 -220
rect 4200 -255 4235 -220
rect 4245 -255 4280 -220
rect 4290 -255 4325 -220
rect 4335 -255 4370 -220
rect 4380 -255 4415 -220
rect 4425 -255 4460 -220
rect 4470 -255 4505 -220
rect 4515 -255 4550 -220
rect 4560 -255 4595 -220
<< mimcap >>
rect 3025 1560 4605 1630
rect 3025 1440 3095 1560
rect 3215 1440 3260 1560
rect 3380 1440 3425 1560
rect 3545 1440 3590 1560
rect 3710 1440 3755 1560
rect 3875 1440 3920 1560
rect 4040 1440 4085 1560
rect 4205 1440 4250 1560
rect 4370 1440 4415 1560
rect 4535 1440 4605 1560
rect 3025 1395 4605 1440
rect 3025 1275 3095 1395
rect 3215 1275 3260 1395
rect 3380 1275 3425 1395
rect 3545 1275 3590 1395
rect 3710 1275 3755 1395
rect 3875 1275 3920 1395
rect 4040 1275 4085 1395
rect 4205 1275 4250 1395
rect 4370 1275 4415 1395
rect 4535 1275 4605 1395
rect 3025 1230 4605 1275
rect 3025 1110 3095 1230
rect 3215 1110 3260 1230
rect 3380 1110 3425 1230
rect 3545 1110 3590 1230
rect 3710 1110 3755 1230
rect 3875 1110 3920 1230
rect 4040 1110 4085 1230
rect 4205 1110 4250 1230
rect 4370 1110 4415 1230
rect 4535 1110 4605 1230
rect 3025 1065 4605 1110
rect 3025 945 3095 1065
rect 3215 945 3260 1065
rect 3380 945 3425 1065
rect 3545 945 3590 1065
rect 3710 945 3755 1065
rect 3875 945 3920 1065
rect 4040 945 4085 1065
rect 4205 945 4250 1065
rect 4370 945 4415 1065
rect 4535 945 4605 1065
rect 3025 900 4605 945
rect 3025 780 3095 900
rect 3215 780 3260 900
rect 3380 780 3425 900
rect 3545 780 3590 900
rect 3710 780 3755 900
rect 3875 780 3920 900
rect 4040 780 4085 900
rect 4205 780 4250 900
rect 4370 780 4415 900
rect 4535 780 4605 900
rect 3025 735 4605 780
rect 3025 615 3095 735
rect 3215 615 3260 735
rect 3380 615 3425 735
rect 3545 615 3590 735
rect 3710 615 3755 735
rect 3875 615 3920 735
rect 4040 615 4085 735
rect 4205 615 4250 735
rect 4370 615 4415 735
rect 4535 615 4605 735
rect 3025 570 4605 615
rect 3025 450 3095 570
rect 3215 450 3260 570
rect 3380 450 3425 570
rect 3545 450 3590 570
rect 3710 450 3755 570
rect 3875 450 3920 570
rect 4040 450 4085 570
rect 4205 450 4250 570
rect 4370 450 4415 570
rect 4535 450 4605 570
rect 3025 405 4605 450
rect 3025 285 3095 405
rect 3215 285 3260 405
rect 3380 285 3425 405
rect 3545 285 3590 405
rect 3710 285 3755 405
rect 3875 285 3920 405
rect 4040 285 4085 405
rect 4205 285 4250 405
rect 4370 285 4415 405
rect 4535 285 4605 405
rect 3025 240 4605 285
rect 3025 120 3095 240
rect 3215 120 3260 240
rect 3380 120 3425 240
rect 3545 120 3590 240
rect 3710 120 3755 240
rect 3875 120 3920 240
rect 4040 120 4085 240
rect 4205 120 4250 240
rect 4370 120 4415 240
rect 4535 120 4605 240
rect 3025 50 4605 120
<< mimcapcontact >>
rect 3095 1440 3215 1560
rect 3260 1440 3380 1560
rect 3425 1440 3545 1560
rect 3590 1440 3710 1560
rect 3755 1440 3875 1560
rect 3920 1440 4040 1560
rect 4085 1440 4205 1560
rect 4250 1440 4370 1560
rect 4415 1440 4535 1560
rect 3095 1275 3215 1395
rect 3260 1275 3380 1395
rect 3425 1275 3545 1395
rect 3590 1275 3710 1395
rect 3755 1275 3875 1395
rect 3920 1275 4040 1395
rect 4085 1275 4205 1395
rect 4250 1275 4370 1395
rect 4415 1275 4535 1395
rect 3095 1110 3215 1230
rect 3260 1110 3380 1230
rect 3425 1110 3545 1230
rect 3590 1110 3710 1230
rect 3755 1110 3875 1230
rect 3920 1110 4040 1230
rect 4085 1110 4205 1230
rect 4250 1110 4370 1230
rect 4415 1110 4535 1230
rect 3095 945 3215 1065
rect 3260 945 3380 1065
rect 3425 945 3545 1065
rect 3590 945 3710 1065
rect 3755 945 3875 1065
rect 3920 945 4040 1065
rect 4085 945 4205 1065
rect 4250 945 4370 1065
rect 4415 945 4535 1065
rect 3095 780 3215 900
rect 3260 780 3380 900
rect 3425 780 3545 900
rect 3590 780 3710 900
rect 3755 780 3875 900
rect 3920 780 4040 900
rect 4085 780 4205 900
rect 4250 780 4370 900
rect 4415 780 4535 900
rect 3095 615 3215 735
rect 3260 615 3380 735
rect 3425 615 3545 735
rect 3590 615 3710 735
rect 3755 615 3875 735
rect 3920 615 4040 735
rect 4085 615 4205 735
rect 4250 615 4370 735
rect 4415 615 4535 735
rect 3095 450 3215 570
rect 3260 450 3380 570
rect 3425 450 3545 570
rect 3590 450 3710 570
rect 3755 450 3875 570
rect 3920 450 4040 570
rect 4085 450 4205 570
rect 4250 450 4370 570
rect 4415 450 4535 570
rect 3095 285 3215 405
rect 3260 285 3380 405
rect 3425 285 3545 405
rect 3590 285 3710 405
rect 3755 285 3875 405
rect 3920 285 4040 405
rect 4085 285 4205 405
rect 4250 285 4370 405
rect 4415 285 4535 405
rect 3095 120 3215 240
rect 3260 120 3380 240
rect 3425 120 3545 240
rect 3590 120 3710 240
rect 3755 120 3875 240
rect 3920 120 4040 240
rect 4085 120 4205 240
rect 4250 120 4370 240
rect 4415 120 4535 240
<< metal4 >>
rect 2770 1640 4620 1645
rect 2770 1605 2780 1640
rect 2815 1605 2830 1640
rect 2865 1605 2880 1640
rect 2915 1605 2930 1640
rect 2965 1605 4620 1640
rect 2770 1600 4620 1605
rect 3010 1560 4620 1600
rect 3010 1440 3095 1560
rect 3215 1440 3260 1560
rect 3380 1440 3425 1560
rect 3545 1440 3590 1560
rect 3710 1440 3755 1560
rect 3875 1440 3920 1560
rect 4040 1440 4085 1560
rect 4205 1440 4250 1560
rect 4370 1440 4415 1560
rect 4535 1440 4620 1560
rect 3010 1395 4620 1440
rect 3010 1275 3095 1395
rect 3215 1275 3260 1395
rect 3380 1275 3425 1395
rect 3545 1275 3590 1395
rect 3710 1275 3755 1395
rect 3875 1275 3920 1395
rect 4040 1275 4085 1395
rect 4205 1275 4250 1395
rect 4370 1275 4415 1395
rect 4535 1275 4620 1395
rect 3010 1230 4620 1275
rect 3010 1110 3095 1230
rect 3215 1110 3260 1230
rect 3380 1110 3425 1230
rect 3545 1110 3590 1230
rect 3710 1110 3755 1230
rect 3875 1110 3920 1230
rect 4040 1110 4085 1230
rect 4205 1110 4250 1230
rect 4370 1110 4415 1230
rect 4535 1110 4620 1230
rect 3010 1065 4620 1110
rect 3010 945 3095 1065
rect 3215 945 3260 1065
rect 3380 945 3425 1065
rect 3545 945 3590 1065
rect 3710 945 3755 1065
rect 3875 945 3920 1065
rect 4040 945 4085 1065
rect 4205 945 4250 1065
rect 4370 945 4415 1065
rect 4535 945 4620 1065
rect 3010 900 4620 945
rect 3010 780 3095 900
rect 3215 780 3260 900
rect 3380 780 3425 900
rect 3545 780 3590 900
rect 3710 780 3755 900
rect 3875 780 3920 900
rect 4040 780 4085 900
rect 4205 780 4250 900
rect 4370 780 4415 900
rect 4535 780 4620 900
rect 3010 735 4620 780
rect 3010 615 3095 735
rect 3215 615 3260 735
rect 3380 615 3425 735
rect 3545 615 3590 735
rect 3710 615 3755 735
rect 3875 615 3920 735
rect 4040 615 4085 735
rect 4205 615 4250 735
rect 4370 615 4415 735
rect 4535 615 4620 735
rect 3010 570 4620 615
rect 3010 450 3095 570
rect 3215 450 3260 570
rect 3380 450 3425 570
rect 3545 450 3590 570
rect 3710 450 3755 570
rect 3875 450 3920 570
rect 4040 450 4085 570
rect 4205 450 4250 570
rect 4370 450 4415 570
rect 4535 450 4620 570
rect 3010 405 4620 450
rect 3010 285 3095 405
rect 3215 285 3260 405
rect 3380 285 3425 405
rect 3545 285 3590 405
rect 3710 285 3755 405
rect 3875 285 3920 405
rect 4040 285 4085 405
rect 4205 285 4250 405
rect 4370 285 4415 405
rect 4535 285 4620 405
rect 3010 240 4620 285
rect 3010 120 3095 240
rect 3215 120 3260 240
rect 3380 120 3425 240
rect 3545 120 3590 240
rect 3710 120 3755 240
rect 3875 120 3920 240
rect 4040 120 4085 240
rect 4205 120 4250 240
rect 4370 120 4415 240
rect 4535 120 4620 240
rect 3010 35 4620 120
rect 3010 -130 4620 -125
rect 3010 -150 3030 -130
rect 3065 -150 3075 -130
rect 3110 -150 3120 -130
rect 3010 -270 3025 -150
rect 3155 -165 3165 -130
rect 3200 -150 3210 -130
rect 3245 -150 3255 -130
rect 3290 -150 3300 -130
rect 3335 -165 3345 -130
rect 3380 -150 3390 -130
rect 3425 -150 3435 -130
rect 3470 -150 3480 -130
rect 3475 -165 3480 -150
rect 3515 -150 3525 -130
rect 3560 -150 3570 -130
rect 3605 -150 3615 -130
rect 3515 -165 3520 -150
rect 3650 -165 3660 -130
rect 3695 -150 3705 -130
rect 3740 -150 3750 -130
rect 3785 -150 3795 -130
rect 3830 -165 3840 -130
rect 3875 -150 3885 -130
rect 3920 -150 3930 -130
rect 3965 -150 3975 -130
rect 3970 -165 3975 -150
rect 4010 -150 4020 -130
rect 4055 -150 4065 -130
rect 4100 -150 4110 -130
rect 4010 -165 4015 -150
rect 4145 -165 4155 -130
rect 4190 -150 4200 -130
rect 4235 -150 4245 -130
rect 4280 -150 4290 -130
rect 4325 -165 4335 -130
rect 4370 -150 4380 -130
rect 4415 -150 4425 -130
rect 4460 -150 4470 -130
rect 4465 -165 4470 -150
rect 4505 -165 4515 -130
rect 4550 -165 4560 -130
rect 4595 -165 4620 -130
rect 3145 -175 3190 -165
rect 3310 -175 3355 -165
rect 3475 -175 3520 -165
rect 3640 -175 3685 -165
rect 3805 -175 3850 -165
rect 3970 -175 4015 -165
rect 4135 -175 4180 -165
rect 4300 -175 4345 -165
rect 4465 -175 4620 -165
rect 3155 -210 3165 -175
rect 3335 -210 3345 -175
rect 3475 -210 3480 -175
rect 3515 -210 3520 -175
rect 3650 -210 3660 -175
rect 3830 -210 3840 -175
rect 3970 -210 3975 -175
rect 4010 -210 4015 -175
rect 4145 -210 4155 -175
rect 4325 -210 4335 -175
rect 4465 -210 4470 -175
rect 4505 -210 4515 -175
rect 4550 -210 4560 -175
rect 4595 -210 4620 -175
rect 3145 -220 3190 -210
rect 3310 -220 3355 -210
rect 3475 -220 3520 -210
rect 3640 -220 3685 -210
rect 3805 -220 3850 -210
rect 3970 -220 4015 -210
rect 4135 -220 4180 -210
rect 4300 -220 4345 -210
rect 4465 -220 4620 -210
rect 3155 -255 3165 -220
rect 3335 -255 3345 -220
rect 3475 -255 3480 -220
rect 3515 -255 3520 -220
rect 3650 -255 3660 -220
rect 3830 -255 3840 -220
rect 3970 -255 3975 -220
rect 4010 -255 4015 -220
rect 4145 -255 4155 -220
rect 4325 -255 4335 -220
rect 4465 -255 4470 -220
rect 4505 -255 4515 -220
rect 4550 -255 4560 -220
rect 4595 -255 4620 -220
rect 3145 -270 3190 -255
rect 3310 -270 3355 -255
rect 3475 -270 3520 -255
rect 3640 -270 3685 -255
rect 3805 -270 3850 -255
rect 3970 -270 4015 -255
rect 4135 -270 4180 -255
rect 4300 -270 4345 -255
rect 4465 -270 4620 -255
rect 3010 -285 4620 -270
<< via4 >>
rect 3025 -165 3030 -150
rect 3030 -165 3065 -150
rect 3065 -165 3075 -150
rect 3075 -165 3110 -150
rect 3110 -165 3120 -150
rect 3120 -165 3145 -150
rect 3190 -165 3200 -150
rect 3200 -165 3210 -150
rect 3210 -165 3245 -150
rect 3245 -165 3255 -150
rect 3255 -165 3290 -150
rect 3290 -165 3300 -150
rect 3300 -165 3310 -150
rect 3355 -165 3380 -150
rect 3380 -165 3390 -150
rect 3390 -165 3425 -150
rect 3425 -165 3435 -150
rect 3435 -165 3470 -150
rect 3470 -165 3475 -150
rect 3520 -165 3525 -150
rect 3525 -165 3560 -150
rect 3560 -165 3570 -150
rect 3570 -165 3605 -150
rect 3605 -165 3615 -150
rect 3615 -165 3640 -150
rect 3685 -165 3695 -150
rect 3695 -165 3705 -150
rect 3705 -165 3740 -150
rect 3740 -165 3750 -150
rect 3750 -165 3785 -150
rect 3785 -165 3795 -150
rect 3795 -165 3805 -150
rect 3850 -165 3875 -150
rect 3875 -165 3885 -150
rect 3885 -165 3920 -150
rect 3920 -165 3930 -150
rect 3930 -165 3965 -150
rect 3965 -165 3970 -150
rect 4015 -165 4020 -150
rect 4020 -165 4055 -150
rect 4055 -165 4065 -150
rect 4065 -165 4100 -150
rect 4100 -165 4110 -150
rect 4110 -165 4135 -150
rect 4180 -165 4190 -150
rect 4190 -165 4200 -150
rect 4200 -165 4235 -150
rect 4235 -165 4245 -150
rect 4245 -165 4280 -150
rect 4280 -165 4290 -150
rect 4290 -165 4300 -150
rect 4345 -165 4370 -150
rect 4370 -165 4380 -150
rect 4380 -165 4415 -150
rect 4415 -165 4425 -150
rect 4425 -165 4460 -150
rect 4460 -165 4465 -150
rect 3025 -175 3145 -165
rect 3190 -175 3310 -165
rect 3355 -175 3475 -165
rect 3520 -175 3640 -165
rect 3685 -175 3805 -165
rect 3850 -175 3970 -165
rect 4015 -175 4135 -165
rect 4180 -175 4300 -165
rect 4345 -175 4465 -165
rect 3025 -210 3030 -175
rect 3030 -210 3065 -175
rect 3065 -210 3075 -175
rect 3075 -210 3110 -175
rect 3110 -210 3120 -175
rect 3120 -210 3145 -175
rect 3190 -210 3200 -175
rect 3200 -210 3210 -175
rect 3210 -210 3245 -175
rect 3245 -210 3255 -175
rect 3255 -210 3290 -175
rect 3290 -210 3300 -175
rect 3300 -210 3310 -175
rect 3355 -210 3380 -175
rect 3380 -210 3390 -175
rect 3390 -210 3425 -175
rect 3425 -210 3435 -175
rect 3435 -210 3470 -175
rect 3470 -210 3475 -175
rect 3520 -210 3525 -175
rect 3525 -210 3560 -175
rect 3560 -210 3570 -175
rect 3570 -210 3605 -175
rect 3605 -210 3615 -175
rect 3615 -210 3640 -175
rect 3685 -210 3695 -175
rect 3695 -210 3705 -175
rect 3705 -210 3740 -175
rect 3740 -210 3750 -175
rect 3750 -210 3785 -175
rect 3785 -210 3795 -175
rect 3795 -210 3805 -175
rect 3850 -210 3875 -175
rect 3875 -210 3885 -175
rect 3885 -210 3920 -175
rect 3920 -210 3930 -175
rect 3930 -210 3965 -175
rect 3965 -210 3970 -175
rect 4015 -210 4020 -175
rect 4020 -210 4055 -175
rect 4055 -210 4065 -175
rect 4065 -210 4100 -175
rect 4100 -210 4110 -175
rect 4110 -210 4135 -175
rect 4180 -210 4190 -175
rect 4190 -210 4200 -175
rect 4200 -210 4235 -175
rect 4235 -210 4245 -175
rect 4245 -210 4280 -175
rect 4280 -210 4290 -175
rect 4290 -210 4300 -175
rect 4345 -210 4370 -175
rect 4370 -210 4380 -175
rect 4380 -210 4415 -175
rect 4415 -210 4425 -175
rect 4425 -210 4460 -175
rect 4460 -210 4465 -175
rect 3025 -220 3145 -210
rect 3190 -220 3310 -210
rect 3355 -220 3475 -210
rect 3520 -220 3640 -210
rect 3685 -220 3805 -210
rect 3850 -220 3970 -210
rect 4015 -220 4135 -210
rect 4180 -220 4300 -210
rect 4345 -220 4465 -210
rect 3025 -255 3030 -220
rect 3030 -255 3065 -220
rect 3065 -255 3075 -220
rect 3075 -255 3110 -220
rect 3110 -255 3120 -220
rect 3120 -255 3145 -220
rect 3190 -255 3200 -220
rect 3200 -255 3210 -220
rect 3210 -255 3245 -220
rect 3245 -255 3255 -220
rect 3255 -255 3290 -220
rect 3290 -255 3300 -220
rect 3300 -255 3310 -220
rect 3355 -255 3380 -220
rect 3380 -255 3390 -220
rect 3390 -255 3425 -220
rect 3425 -255 3435 -220
rect 3435 -255 3470 -220
rect 3470 -255 3475 -220
rect 3520 -255 3525 -220
rect 3525 -255 3560 -220
rect 3560 -255 3570 -220
rect 3570 -255 3605 -220
rect 3605 -255 3615 -220
rect 3615 -255 3640 -220
rect 3685 -255 3695 -220
rect 3695 -255 3705 -220
rect 3705 -255 3740 -220
rect 3740 -255 3750 -220
rect 3750 -255 3785 -220
rect 3785 -255 3795 -220
rect 3795 -255 3805 -220
rect 3850 -255 3875 -220
rect 3875 -255 3885 -220
rect 3885 -255 3920 -220
rect 3920 -255 3930 -220
rect 3930 -255 3965 -220
rect 3965 -255 3970 -220
rect 4015 -255 4020 -220
rect 4020 -255 4055 -220
rect 4055 -255 4065 -220
rect 4065 -255 4100 -220
rect 4100 -255 4110 -220
rect 4110 -255 4135 -220
rect 4180 -255 4190 -220
rect 4190 -255 4200 -220
rect 4200 -255 4235 -220
rect 4235 -255 4245 -220
rect 4245 -255 4280 -220
rect 4280 -255 4290 -220
rect 4290 -255 4300 -220
rect 4345 -255 4370 -220
rect 4370 -255 4380 -220
rect 4380 -255 4415 -220
rect 4415 -255 4425 -220
rect 4425 -255 4460 -220
rect 4460 -255 4465 -220
rect 3025 -270 3145 -255
rect 3190 -270 3310 -255
rect 3355 -270 3475 -255
rect 3520 -270 3640 -255
rect 3685 -270 3805 -255
rect 3850 -270 3970 -255
rect 4015 -270 4135 -255
rect 4180 -270 4300 -255
rect 4345 -270 4465 -255
<< mimcap2 >>
rect 3025 1560 4605 1630
rect 3025 1440 3095 1560
rect 3215 1440 3260 1560
rect 3380 1440 3425 1560
rect 3545 1440 3590 1560
rect 3710 1440 3755 1560
rect 3875 1440 3920 1560
rect 4040 1440 4085 1560
rect 4205 1440 4250 1560
rect 4370 1440 4415 1560
rect 4535 1440 4605 1560
rect 3025 1395 4605 1440
rect 3025 1275 3095 1395
rect 3215 1275 3260 1395
rect 3380 1275 3425 1395
rect 3545 1275 3590 1395
rect 3710 1275 3755 1395
rect 3875 1275 3920 1395
rect 4040 1275 4085 1395
rect 4205 1275 4250 1395
rect 4370 1275 4415 1395
rect 4535 1275 4605 1395
rect 3025 1230 4605 1275
rect 3025 1110 3095 1230
rect 3215 1110 3260 1230
rect 3380 1110 3425 1230
rect 3545 1110 3590 1230
rect 3710 1110 3755 1230
rect 3875 1110 3920 1230
rect 4040 1110 4085 1230
rect 4205 1110 4250 1230
rect 4370 1110 4415 1230
rect 4535 1110 4605 1230
rect 3025 1065 4605 1110
rect 3025 945 3095 1065
rect 3215 945 3260 1065
rect 3380 945 3425 1065
rect 3545 945 3590 1065
rect 3710 945 3755 1065
rect 3875 945 3920 1065
rect 4040 945 4085 1065
rect 4205 945 4250 1065
rect 4370 945 4415 1065
rect 4535 945 4605 1065
rect 3025 900 4605 945
rect 3025 780 3095 900
rect 3215 780 3260 900
rect 3380 780 3425 900
rect 3545 780 3590 900
rect 3710 780 3755 900
rect 3875 780 3920 900
rect 4040 780 4085 900
rect 4205 780 4250 900
rect 4370 780 4415 900
rect 4535 780 4605 900
rect 3025 735 4605 780
rect 3025 615 3095 735
rect 3215 615 3260 735
rect 3380 615 3425 735
rect 3545 615 3590 735
rect 3710 615 3755 735
rect 3875 615 3920 735
rect 4040 615 4085 735
rect 4205 615 4250 735
rect 4370 615 4415 735
rect 4535 615 4605 735
rect 3025 570 4605 615
rect 3025 450 3095 570
rect 3215 450 3260 570
rect 3380 450 3425 570
rect 3545 450 3590 570
rect 3710 450 3755 570
rect 3875 450 3920 570
rect 4040 450 4085 570
rect 4205 450 4250 570
rect 4370 450 4415 570
rect 4535 450 4605 570
rect 3025 405 4605 450
rect 3025 285 3095 405
rect 3215 285 3260 405
rect 3380 285 3425 405
rect 3545 285 3590 405
rect 3710 285 3755 405
rect 3875 285 3920 405
rect 4040 285 4085 405
rect 4205 285 4250 405
rect 4370 285 4415 405
rect 4535 285 4605 405
rect 3025 240 4605 285
rect 3025 120 3095 240
rect 3215 120 3260 240
rect 3380 120 3425 240
rect 3545 120 3590 240
rect 3710 120 3755 240
rect 3875 120 3920 240
rect 4040 120 4085 240
rect 4205 120 4250 240
rect 4370 120 4415 240
rect 4535 120 4605 240
rect 3025 50 4605 120
<< mimcap2contact >>
rect 3095 1440 3215 1560
rect 3260 1440 3380 1560
rect 3425 1440 3545 1560
rect 3590 1440 3710 1560
rect 3755 1440 3875 1560
rect 3920 1440 4040 1560
rect 4085 1440 4205 1560
rect 4250 1440 4370 1560
rect 4415 1440 4535 1560
rect 3095 1275 3215 1395
rect 3260 1275 3380 1395
rect 3425 1275 3545 1395
rect 3590 1275 3710 1395
rect 3755 1275 3875 1395
rect 3920 1275 4040 1395
rect 4085 1275 4205 1395
rect 4250 1275 4370 1395
rect 4415 1275 4535 1395
rect 3095 1110 3215 1230
rect 3260 1110 3380 1230
rect 3425 1110 3545 1230
rect 3590 1110 3710 1230
rect 3755 1110 3875 1230
rect 3920 1110 4040 1230
rect 4085 1110 4205 1230
rect 4250 1110 4370 1230
rect 4415 1110 4535 1230
rect 3095 945 3215 1065
rect 3260 945 3380 1065
rect 3425 945 3545 1065
rect 3590 945 3710 1065
rect 3755 945 3875 1065
rect 3920 945 4040 1065
rect 4085 945 4205 1065
rect 4250 945 4370 1065
rect 4415 945 4535 1065
rect 3095 780 3215 900
rect 3260 780 3380 900
rect 3425 780 3545 900
rect 3590 780 3710 900
rect 3755 780 3875 900
rect 3920 780 4040 900
rect 4085 780 4205 900
rect 4250 780 4370 900
rect 4415 780 4535 900
rect 3095 615 3215 735
rect 3260 615 3380 735
rect 3425 615 3545 735
rect 3590 615 3710 735
rect 3755 615 3875 735
rect 3920 615 4040 735
rect 4085 615 4205 735
rect 4250 615 4370 735
rect 4415 615 4535 735
rect 3095 450 3215 570
rect 3260 450 3380 570
rect 3425 450 3545 570
rect 3590 450 3710 570
rect 3755 450 3875 570
rect 3920 450 4040 570
rect 4085 450 4205 570
rect 4250 450 4370 570
rect 4415 450 4535 570
rect 3095 285 3215 405
rect 3260 285 3380 405
rect 3425 285 3545 405
rect 3590 285 3710 405
rect 3755 285 3875 405
rect 3920 285 4040 405
rect 4085 285 4205 405
rect 4250 285 4370 405
rect 4415 285 4535 405
rect 3095 120 3215 240
rect 3260 120 3380 240
rect 3425 120 3545 240
rect 3590 120 3710 240
rect 3755 120 3875 240
rect 3920 120 4040 240
rect 4085 120 4205 240
rect 4250 120 4370 240
rect 4415 120 4535 240
<< metal5 >>
rect 3010 1560 4620 1645
rect 3010 1440 3095 1560
rect 3215 1440 3260 1560
rect 3380 1440 3425 1560
rect 3545 1440 3590 1560
rect 3710 1440 3755 1560
rect 3875 1440 3920 1560
rect 4040 1440 4085 1560
rect 4205 1440 4250 1560
rect 4370 1440 4415 1560
rect 4535 1440 4620 1560
rect 3010 1395 4620 1440
rect 3010 1275 3095 1395
rect 3215 1275 3260 1395
rect 3380 1275 3425 1395
rect 3545 1275 3590 1395
rect 3710 1275 3755 1395
rect 3875 1275 3920 1395
rect 4040 1275 4085 1395
rect 4205 1275 4250 1395
rect 4370 1275 4415 1395
rect 4535 1275 4620 1395
rect 3010 1230 4620 1275
rect 3010 1110 3095 1230
rect 3215 1110 3260 1230
rect 3380 1110 3425 1230
rect 3545 1110 3590 1230
rect 3710 1110 3755 1230
rect 3875 1110 3920 1230
rect 4040 1110 4085 1230
rect 4205 1110 4250 1230
rect 4370 1110 4415 1230
rect 4535 1110 4620 1230
rect 3010 1065 4620 1110
rect 3010 945 3095 1065
rect 3215 945 3260 1065
rect 3380 945 3425 1065
rect 3545 945 3590 1065
rect 3710 945 3755 1065
rect 3875 945 3920 1065
rect 4040 945 4085 1065
rect 4205 945 4250 1065
rect 4370 945 4415 1065
rect 4535 945 4620 1065
rect 3010 900 4620 945
rect 3010 780 3095 900
rect 3215 780 3260 900
rect 3380 780 3425 900
rect 3545 780 3590 900
rect 3710 780 3755 900
rect 3875 780 3920 900
rect 4040 780 4085 900
rect 4205 780 4250 900
rect 4370 780 4415 900
rect 4535 780 4620 900
rect 3010 735 4620 780
rect 3010 615 3095 735
rect 3215 615 3260 735
rect 3380 615 3425 735
rect 3545 615 3590 735
rect 3710 615 3755 735
rect 3875 615 3920 735
rect 4040 615 4085 735
rect 4205 615 4250 735
rect 4370 615 4415 735
rect 4535 615 4620 735
rect 3010 570 4620 615
rect 3010 450 3095 570
rect 3215 450 3260 570
rect 3380 450 3425 570
rect 3545 450 3590 570
rect 3710 450 3755 570
rect 3875 450 3920 570
rect 4040 450 4085 570
rect 4205 450 4250 570
rect 4370 450 4415 570
rect 4535 450 4620 570
rect 3010 405 4620 450
rect 3010 285 3095 405
rect 3215 285 3260 405
rect 3380 285 3425 405
rect 3545 285 3590 405
rect 3710 285 3755 405
rect 3875 285 3920 405
rect 4040 285 4085 405
rect 4205 285 4250 405
rect 4370 285 4415 405
rect 4535 285 4620 405
rect 3010 240 4620 285
rect 3010 120 3095 240
rect 3215 120 3260 240
rect 3380 120 3425 240
rect 3545 120 3590 240
rect 3710 120 3755 240
rect 3875 120 3920 240
rect 4040 120 4085 240
rect 4205 120 4250 240
rect 4370 120 4415 240
rect 4535 120 4620 240
rect 3010 -150 4620 120
rect 3010 -270 3025 -150
rect 3145 -270 3190 -150
rect 3310 -270 3355 -150
rect 3475 -270 3520 -150
rect 3640 -270 3685 -150
rect 3805 -270 3850 -150
rect 3970 -270 4015 -150
rect 4135 -270 4180 -150
rect 4300 -270 4345 -150
rect 4465 -270 4620 -150
rect 3010 -285 4620 -270
<< labels >>
rlabel metal5 3825 -280 3825 -280 1 GND
port 2 n
rlabel metal1 665 280 665 280 1 GND
port 2 n
rlabel metal4 2990 1640 2990 1640 1 Vb3
port 5 n
rlabel viali 880 125 880 125 1 Vb3_
port 6 n
rlabel metal1 575 15 575 15 1 GND
port 2 n
<< end >>
