magic
tech sky130A
timestamp 1634762988
<< nmos >>
rect 105 -130 2605 -85
rect 105 -225 2605 -180
rect 105 -320 2605 -275
rect 105 -415 2605 -370
rect 105 -510 2605 -465
rect 105 -605 2605 -560
rect 105 -700 2605 -655
rect 105 -795 2605 -750
rect 105 -890 2605 -845
rect 105 -985 2605 -940
rect 105 -1080 2605 -1035
rect 105 -1175 2605 -1130
rect 105 -1270 2605 -1225
rect 105 -1365 2605 -1320
rect 105 -1460 2605 -1415
rect 105 -1555 2605 -1510
rect 105 -1650 2605 -1605
rect 105 -1745 2605 -1700
rect 105 -1840 2605 -1795
rect 105 -1935 2605 -1890
rect 105 -2030 2605 -1985
rect 105 -2125 2605 -2080
rect 105 -2220 2605 -2175
rect 105 -2315 2605 -2270
rect 105 -2410 2605 -2365
rect 105 -2505 2605 -2460
<< nmoslvt >>
rect 175 2230 2675 2262
rect 175 2148 2675 2180
rect 175 2066 2675 2098
rect 175 1984 2675 2016
rect 175 1902 2675 1934
rect 175 1820 2675 1852
rect 175 1738 2675 1770
rect 175 1656 2675 1688
rect 175 1574 2675 1606
rect 175 1492 2675 1524
rect 175 1410 2675 1442
rect 175 1328 2675 1360
rect 175 1246 2675 1278
rect 175 1164 2675 1196
rect 175 1082 2675 1114
rect 175 1000 2675 1032
rect 175 918 2675 950
rect 175 836 2675 868
rect 175 754 2675 786
rect 175 672 2675 704
rect 175 590 2675 622
rect 175 508 2675 540
rect 175 426 2675 458
rect 175 344 2675 376
rect 175 262 2675 294
rect 175 180 2675 212
<< ndiff >>
rect 175 2297 2675 2307
rect 175 2277 200 2297
rect 220 2277 240 2297
rect 260 2277 280 2297
rect 300 2277 320 2297
rect 340 2277 360 2297
rect 380 2277 400 2297
rect 420 2277 440 2297
rect 460 2277 480 2297
rect 500 2277 520 2297
rect 540 2277 560 2297
rect 580 2277 600 2297
rect 620 2277 640 2297
rect 660 2277 680 2297
rect 700 2277 720 2297
rect 740 2277 760 2297
rect 780 2277 800 2297
rect 820 2277 840 2297
rect 860 2277 880 2297
rect 900 2277 920 2297
rect 940 2277 960 2297
rect 980 2277 1000 2297
rect 1020 2277 1040 2297
rect 1060 2277 1080 2297
rect 1100 2277 1120 2297
rect 1140 2277 1160 2297
rect 1180 2277 1200 2297
rect 1220 2277 1240 2297
rect 1260 2277 1280 2297
rect 1300 2277 1320 2297
rect 1340 2277 1360 2297
rect 1380 2277 1400 2297
rect 1420 2277 1440 2297
rect 1460 2277 1480 2297
rect 1500 2277 1520 2297
rect 1540 2277 1560 2297
rect 1580 2277 1600 2297
rect 1620 2277 1640 2297
rect 1660 2277 1680 2297
rect 1700 2277 1720 2297
rect 1740 2277 1760 2297
rect 1780 2277 1800 2297
rect 1820 2277 1840 2297
rect 1860 2277 1880 2297
rect 1900 2277 1920 2297
rect 1940 2277 1960 2297
rect 1980 2277 2000 2297
rect 2020 2277 2040 2297
rect 2060 2277 2080 2297
rect 2100 2277 2120 2297
rect 2140 2277 2160 2297
rect 2180 2277 2200 2297
rect 2220 2277 2240 2297
rect 2260 2277 2280 2297
rect 2300 2277 2320 2297
rect 2340 2277 2360 2297
rect 2380 2277 2400 2297
rect 2420 2277 2440 2297
rect 2460 2277 2480 2297
rect 2500 2277 2520 2297
rect 2540 2277 2560 2297
rect 2580 2277 2600 2297
rect 2620 2277 2640 2297
rect 2660 2277 2675 2297
rect 175 2262 2675 2277
rect 175 2215 2675 2230
rect 175 2195 200 2215
rect 220 2195 240 2215
rect 260 2195 280 2215
rect 300 2195 320 2215
rect 340 2195 360 2215
rect 380 2195 400 2215
rect 420 2195 440 2215
rect 460 2195 480 2215
rect 500 2195 520 2215
rect 540 2195 560 2215
rect 580 2195 600 2215
rect 620 2195 640 2215
rect 660 2195 680 2215
rect 700 2195 720 2215
rect 740 2195 760 2215
rect 780 2195 800 2215
rect 820 2195 840 2215
rect 860 2195 880 2215
rect 900 2195 920 2215
rect 940 2195 960 2215
rect 980 2195 1000 2215
rect 1020 2195 1040 2215
rect 1060 2195 1080 2215
rect 1100 2195 1120 2215
rect 1140 2195 1160 2215
rect 1180 2195 1200 2215
rect 1220 2195 1240 2215
rect 1260 2195 1280 2215
rect 1300 2195 1320 2215
rect 1340 2195 1360 2215
rect 1380 2195 1400 2215
rect 1420 2195 1440 2215
rect 1460 2195 1480 2215
rect 1500 2195 1520 2215
rect 1540 2195 1560 2215
rect 1580 2195 1600 2215
rect 1620 2195 1640 2215
rect 1660 2195 1680 2215
rect 1700 2195 1720 2215
rect 1740 2195 1760 2215
rect 1780 2195 1800 2215
rect 1820 2195 1840 2215
rect 1860 2195 1880 2215
rect 1900 2195 1920 2215
rect 1940 2195 1960 2215
rect 1980 2195 2000 2215
rect 2020 2195 2040 2215
rect 2060 2195 2080 2215
rect 2100 2195 2120 2215
rect 2140 2195 2160 2215
rect 2180 2195 2200 2215
rect 2220 2195 2240 2215
rect 2260 2195 2280 2215
rect 2300 2195 2320 2215
rect 2340 2195 2360 2215
rect 2380 2195 2400 2215
rect 2420 2195 2440 2215
rect 2460 2195 2480 2215
rect 2500 2195 2520 2215
rect 2540 2195 2560 2215
rect 2580 2195 2600 2215
rect 2620 2195 2640 2215
rect 2660 2195 2675 2215
rect 175 2180 2675 2195
rect 175 2133 2675 2148
rect 175 2113 200 2133
rect 220 2113 240 2133
rect 260 2113 280 2133
rect 300 2113 320 2133
rect 340 2113 360 2133
rect 380 2113 400 2133
rect 420 2113 440 2133
rect 460 2113 480 2133
rect 500 2113 520 2133
rect 540 2113 560 2133
rect 580 2113 600 2133
rect 620 2113 640 2133
rect 660 2113 680 2133
rect 700 2113 720 2133
rect 740 2113 760 2133
rect 780 2113 800 2133
rect 820 2113 840 2133
rect 860 2113 880 2133
rect 900 2113 920 2133
rect 940 2113 960 2133
rect 980 2113 1000 2133
rect 1020 2113 1040 2133
rect 1060 2113 1080 2133
rect 1100 2113 1120 2133
rect 1140 2113 1160 2133
rect 1180 2113 1200 2133
rect 1220 2113 1240 2133
rect 1260 2113 1280 2133
rect 1300 2113 1320 2133
rect 1340 2113 1360 2133
rect 1380 2113 1400 2133
rect 1420 2113 1440 2133
rect 1460 2113 1480 2133
rect 1500 2113 1520 2133
rect 1540 2113 1560 2133
rect 1580 2113 1600 2133
rect 1620 2113 1640 2133
rect 1660 2113 1680 2133
rect 1700 2113 1720 2133
rect 1740 2113 1760 2133
rect 1780 2113 1800 2133
rect 1820 2113 1840 2133
rect 1860 2113 1880 2133
rect 1900 2113 1920 2133
rect 1940 2113 1960 2133
rect 1980 2113 2000 2133
rect 2020 2113 2040 2133
rect 2060 2113 2080 2133
rect 2100 2113 2120 2133
rect 2140 2113 2160 2133
rect 2180 2113 2200 2133
rect 2220 2113 2240 2133
rect 2260 2113 2280 2133
rect 2300 2113 2320 2133
rect 2340 2113 2360 2133
rect 2380 2113 2400 2133
rect 2420 2113 2440 2133
rect 2460 2113 2480 2133
rect 2500 2113 2520 2133
rect 2540 2113 2560 2133
rect 2580 2113 2600 2133
rect 2620 2113 2640 2133
rect 2660 2113 2675 2133
rect 175 2098 2675 2113
rect 175 2051 2675 2066
rect 175 2031 200 2051
rect 220 2031 240 2051
rect 260 2031 280 2051
rect 300 2031 320 2051
rect 340 2031 360 2051
rect 380 2031 400 2051
rect 420 2031 440 2051
rect 460 2031 480 2051
rect 500 2031 520 2051
rect 540 2031 560 2051
rect 580 2031 600 2051
rect 620 2031 640 2051
rect 660 2031 680 2051
rect 700 2031 720 2051
rect 740 2031 760 2051
rect 780 2031 800 2051
rect 820 2031 840 2051
rect 860 2031 880 2051
rect 900 2031 920 2051
rect 940 2031 960 2051
rect 980 2031 1000 2051
rect 1020 2031 1040 2051
rect 1060 2031 1080 2051
rect 1100 2031 1120 2051
rect 1140 2031 1160 2051
rect 1180 2031 1200 2051
rect 1220 2031 1240 2051
rect 1260 2031 1280 2051
rect 1300 2031 1320 2051
rect 1340 2031 1360 2051
rect 1380 2031 1400 2051
rect 1420 2031 1440 2051
rect 1460 2031 1480 2051
rect 1500 2031 1520 2051
rect 1540 2031 1560 2051
rect 1580 2031 1600 2051
rect 1620 2031 1640 2051
rect 1660 2031 1680 2051
rect 1700 2031 1720 2051
rect 1740 2031 1760 2051
rect 1780 2031 1800 2051
rect 1820 2031 1840 2051
rect 1860 2031 1880 2051
rect 1900 2031 1920 2051
rect 1940 2031 1960 2051
rect 1980 2031 2000 2051
rect 2020 2031 2040 2051
rect 2060 2031 2080 2051
rect 2100 2031 2120 2051
rect 2140 2031 2160 2051
rect 2180 2031 2200 2051
rect 2220 2031 2240 2051
rect 2260 2031 2280 2051
rect 2300 2031 2320 2051
rect 2340 2031 2360 2051
rect 2380 2031 2400 2051
rect 2420 2031 2440 2051
rect 2460 2031 2480 2051
rect 2500 2031 2520 2051
rect 2540 2031 2560 2051
rect 2580 2031 2600 2051
rect 2620 2031 2640 2051
rect 2660 2031 2675 2051
rect 175 2016 2675 2031
rect 175 1969 2675 1984
rect 175 1949 200 1969
rect 220 1949 240 1969
rect 260 1949 280 1969
rect 300 1949 320 1969
rect 340 1949 360 1969
rect 380 1949 400 1969
rect 420 1949 440 1969
rect 460 1949 480 1969
rect 500 1949 520 1969
rect 540 1949 560 1969
rect 580 1949 600 1969
rect 620 1949 640 1969
rect 660 1949 680 1969
rect 700 1949 720 1969
rect 740 1949 760 1969
rect 780 1949 800 1969
rect 820 1949 840 1969
rect 860 1949 880 1969
rect 900 1949 920 1969
rect 940 1949 960 1969
rect 980 1949 1000 1969
rect 1020 1949 1040 1969
rect 1060 1949 1080 1969
rect 1100 1949 1120 1969
rect 1140 1949 1160 1969
rect 1180 1949 1200 1969
rect 1220 1949 1240 1969
rect 1260 1949 1280 1969
rect 1300 1949 1320 1969
rect 1340 1949 1360 1969
rect 1380 1949 1400 1969
rect 1420 1949 1440 1969
rect 1460 1949 1480 1969
rect 1500 1949 1520 1969
rect 1540 1949 1560 1969
rect 1580 1949 1600 1969
rect 1620 1949 1640 1969
rect 1660 1949 1680 1969
rect 1700 1949 1720 1969
rect 1740 1949 1760 1969
rect 1780 1949 1800 1969
rect 1820 1949 1840 1969
rect 1860 1949 1880 1969
rect 1900 1949 1920 1969
rect 1940 1949 1960 1969
rect 1980 1949 2000 1969
rect 2020 1949 2040 1969
rect 2060 1949 2080 1969
rect 2100 1949 2120 1969
rect 2140 1949 2160 1969
rect 2180 1949 2200 1969
rect 2220 1949 2240 1969
rect 2260 1949 2280 1969
rect 2300 1949 2320 1969
rect 2340 1949 2360 1969
rect 2380 1949 2400 1969
rect 2420 1949 2440 1969
rect 2460 1949 2480 1969
rect 2500 1949 2520 1969
rect 2540 1949 2560 1969
rect 2580 1949 2600 1969
rect 2620 1949 2640 1969
rect 2660 1949 2675 1969
rect 175 1934 2675 1949
rect 175 1887 2675 1902
rect 175 1867 200 1887
rect 220 1867 240 1887
rect 260 1867 280 1887
rect 300 1867 320 1887
rect 340 1867 360 1887
rect 380 1867 400 1887
rect 420 1867 440 1887
rect 460 1867 480 1887
rect 500 1867 520 1887
rect 540 1867 560 1887
rect 580 1867 600 1887
rect 620 1867 640 1887
rect 660 1867 680 1887
rect 700 1867 720 1887
rect 740 1867 760 1887
rect 780 1867 800 1887
rect 820 1867 840 1887
rect 860 1867 880 1887
rect 900 1867 920 1887
rect 940 1867 960 1887
rect 980 1867 1000 1887
rect 1020 1867 1040 1887
rect 1060 1867 1080 1887
rect 1100 1867 1120 1887
rect 1140 1867 1160 1887
rect 1180 1867 1200 1887
rect 1220 1867 1240 1887
rect 1260 1867 1280 1887
rect 1300 1867 1320 1887
rect 1340 1867 1360 1887
rect 1380 1867 1400 1887
rect 1420 1867 1440 1887
rect 1460 1867 1480 1887
rect 1500 1867 1520 1887
rect 1540 1867 1560 1887
rect 1580 1867 1600 1887
rect 1620 1867 1640 1887
rect 1660 1867 1680 1887
rect 1700 1867 1720 1887
rect 1740 1867 1760 1887
rect 1780 1867 1800 1887
rect 1820 1867 1840 1887
rect 1860 1867 1880 1887
rect 1900 1867 1920 1887
rect 1940 1867 1960 1887
rect 1980 1867 2000 1887
rect 2020 1867 2040 1887
rect 2060 1867 2080 1887
rect 2100 1867 2120 1887
rect 2140 1867 2160 1887
rect 2180 1867 2200 1887
rect 2220 1867 2240 1887
rect 2260 1867 2280 1887
rect 2300 1867 2320 1887
rect 2340 1867 2360 1887
rect 2380 1867 2400 1887
rect 2420 1867 2440 1887
rect 2460 1867 2480 1887
rect 2500 1867 2520 1887
rect 2540 1867 2560 1887
rect 2580 1867 2600 1887
rect 2620 1867 2640 1887
rect 2660 1867 2675 1887
rect 175 1852 2675 1867
rect 175 1805 2675 1820
rect 175 1785 200 1805
rect 220 1785 240 1805
rect 260 1785 280 1805
rect 300 1785 320 1805
rect 340 1785 360 1805
rect 380 1785 400 1805
rect 420 1785 440 1805
rect 460 1785 480 1805
rect 500 1785 520 1805
rect 540 1785 560 1805
rect 580 1785 600 1805
rect 620 1785 640 1805
rect 660 1785 680 1805
rect 700 1785 720 1805
rect 740 1785 760 1805
rect 780 1785 800 1805
rect 820 1785 840 1805
rect 860 1785 880 1805
rect 900 1785 920 1805
rect 940 1785 960 1805
rect 980 1785 1000 1805
rect 1020 1785 1040 1805
rect 1060 1785 1080 1805
rect 1100 1785 1120 1805
rect 1140 1785 1160 1805
rect 1180 1785 1200 1805
rect 1220 1785 1240 1805
rect 1260 1785 1280 1805
rect 1300 1785 1320 1805
rect 1340 1785 1360 1805
rect 1380 1785 1400 1805
rect 1420 1785 1440 1805
rect 1460 1785 1480 1805
rect 1500 1785 1520 1805
rect 1540 1785 1560 1805
rect 1580 1785 1600 1805
rect 1620 1785 1640 1805
rect 1660 1785 1680 1805
rect 1700 1785 1720 1805
rect 1740 1785 1760 1805
rect 1780 1785 1800 1805
rect 1820 1785 1840 1805
rect 1860 1785 1880 1805
rect 1900 1785 1920 1805
rect 1940 1785 1960 1805
rect 1980 1785 2000 1805
rect 2020 1785 2040 1805
rect 2060 1785 2080 1805
rect 2100 1785 2120 1805
rect 2140 1785 2160 1805
rect 2180 1785 2200 1805
rect 2220 1785 2240 1805
rect 2260 1785 2280 1805
rect 2300 1785 2320 1805
rect 2340 1785 2360 1805
rect 2380 1785 2400 1805
rect 2420 1785 2440 1805
rect 2460 1785 2480 1805
rect 2500 1785 2520 1805
rect 2540 1785 2560 1805
rect 2580 1785 2600 1805
rect 2620 1785 2640 1805
rect 2660 1785 2675 1805
rect 175 1770 2675 1785
rect 175 1723 2675 1738
rect 175 1703 200 1723
rect 220 1703 240 1723
rect 260 1703 280 1723
rect 300 1703 320 1723
rect 340 1703 360 1723
rect 380 1703 400 1723
rect 420 1703 440 1723
rect 460 1703 480 1723
rect 500 1703 520 1723
rect 540 1703 560 1723
rect 580 1703 600 1723
rect 620 1703 640 1723
rect 660 1703 680 1723
rect 700 1703 720 1723
rect 740 1703 760 1723
rect 780 1703 800 1723
rect 820 1703 840 1723
rect 860 1703 880 1723
rect 900 1703 920 1723
rect 940 1703 960 1723
rect 980 1703 1000 1723
rect 1020 1703 1040 1723
rect 1060 1703 1080 1723
rect 1100 1703 1120 1723
rect 1140 1703 1160 1723
rect 1180 1703 1200 1723
rect 1220 1703 1240 1723
rect 1260 1703 1280 1723
rect 1300 1703 1320 1723
rect 1340 1703 1360 1723
rect 1380 1703 1400 1723
rect 1420 1703 1440 1723
rect 1460 1703 1480 1723
rect 1500 1703 1520 1723
rect 1540 1703 1560 1723
rect 1580 1703 1600 1723
rect 1620 1703 1640 1723
rect 1660 1703 1680 1723
rect 1700 1703 1720 1723
rect 1740 1703 1760 1723
rect 1780 1703 1800 1723
rect 1820 1703 1840 1723
rect 1860 1703 1880 1723
rect 1900 1703 1920 1723
rect 1940 1703 1960 1723
rect 1980 1703 2000 1723
rect 2020 1703 2040 1723
rect 2060 1703 2080 1723
rect 2100 1703 2120 1723
rect 2140 1703 2160 1723
rect 2180 1703 2200 1723
rect 2220 1703 2240 1723
rect 2260 1703 2280 1723
rect 2300 1703 2320 1723
rect 2340 1703 2360 1723
rect 2380 1703 2400 1723
rect 2420 1703 2440 1723
rect 2460 1703 2480 1723
rect 2500 1703 2520 1723
rect 2540 1703 2560 1723
rect 2580 1703 2600 1723
rect 2620 1703 2640 1723
rect 2660 1703 2675 1723
rect 175 1688 2675 1703
rect 175 1641 2675 1656
rect 175 1621 200 1641
rect 220 1621 240 1641
rect 260 1621 280 1641
rect 300 1621 320 1641
rect 340 1621 360 1641
rect 380 1621 400 1641
rect 420 1621 440 1641
rect 460 1621 480 1641
rect 500 1621 520 1641
rect 540 1621 560 1641
rect 580 1621 600 1641
rect 620 1621 640 1641
rect 660 1621 680 1641
rect 700 1621 720 1641
rect 740 1621 760 1641
rect 780 1621 800 1641
rect 820 1621 840 1641
rect 860 1621 880 1641
rect 900 1621 920 1641
rect 940 1621 960 1641
rect 980 1621 1000 1641
rect 1020 1621 1040 1641
rect 1060 1621 1080 1641
rect 1100 1621 1120 1641
rect 1140 1621 1160 1641
rect 1180 1621 1200 1641
rect 1220 1621 1240 1641
rect 1260 1621 1280 1641
rect 1300 1621 1320 1641
rect 1340 1621 1360 1641
rect 1380 1621 1400 1641
rect 1420 1621 1440 1641
rect 1460 1621 1480 1641
rect 1500 1621 1520 1641
rect 1540 1621 1560 1641
rect 1580 1621 1600 1641
rect 1620 1621 1640 1641
rect 1660 1621 1680 1641
rect 1700 1621 1720 1641
rect 1740 1621 1760 1641
rect 1780 1621 1800 1641
rect 1820 1621 1840 1641
rect 1860 1621 1880 1641
rect 1900 1621 1920 1641
rect 1940 1621 1960 1641
rect 1980 1621 2000 1641
rect 2020 1621 2040 1641
rect 2060 1621 2080 1641
rect 2100 1621 2120 1641
rect 2140 1621 2160 1641
rect 2180 1621 2200 1641
rect 2220 1621 2240 1641
rect 2260 1621 2280 1641
rect 2300 1621 2320 1641
rect 2340 1621 2360 1641
rect 2380 1621 2400 1641
rect 2420 1621 2440 1641
rect 2460 1621 2480 1641
rect 2500 1621 2520 1641
rect 2540 1621 2560 1641
rect 2580 1621 2600 1641
rect 2620 1621 2640 1641
rect 2660 1621 2675 1641
rect 175 1606 2675 1621
rect 175 1559 2675 1574
rect 175 1539 200 1559
rect 220 1539 240 1559
rect 260 1539 280 1559
rect 300 1539 320 1559
rect 340 1539 360 1559
rect 380 1539 400 1559
rect 420 1539 440 1559
rect 460 1539 480 1559
rect 500 1539 520 1559
rect 540 1539 560 1559
rect 580 1539 600 1559
rect 620 1539 640 1559
rect 660 1539 680 1559
rect 700 1539 720 1559
rect 740 1539 760 1559
rect 780 1539 800 1559
rect 820 1539 840 1559
rect 860 1539 880 1559
rect 900 1539 920 1559
rect 940 1539 960 1559
rect 980 1539 1000 1559
rect 1020 1539 1040 1559
rect 1060 1539 1080 1559
rect 1100 1539 1120 1559
rect 1140 1539 1160 1559
rect 1180 1539 1200 1559
rect 1220 1539 1240 1559
rect 1260 1539 1280 1559
rect 1300 1539 1320 1559
rect 1340 1539 1360 1559
rect 1380 1539 1400 1559
rect 1420 1539 1440 1559
rect 1460 1539 1480 1559
rect 1500 1539 1520 1559
rect 1540 1539 1560 1559
rect 1580 1539 1600 1559
rect 1620 1539 1640 1559
rect 1660 1539 1680 1559
rect 1700 1539 1720 1559
rect 1740 1539 1760 1559
rect 1780 1539 1800 1559
rect 1820 1539 1840 1559
rect 1860 1539 1880 1559
rect 1900 1539 1920 1559
rect 1940 1539 1960 1559
rect 1980 1539 2000 1559
rect 2020 1539 2040 1559
rect 2060 1539 2080 1559
rect 2100 1539 2120 1559
rect 2140 1539 2160 1559
rect 2180 1539 2200 1559
rect 2220 1539 2240 1559
rect 2260 1539 2280 1559
rect 2300 1539 2320 1559
rect 2340 1539 2360 1559
rect 2380 1539 2400 1559
rect 2420 1539 2440 1559
rect 2460 1539 2480 1559
rect 2500 1539 2520 1559
rect 2540 1539 2560 1559
rect 2580 1539 2600 1559
rect 2620 1539 2640 1559
rect 2660 1539 2675 1559
rect 175 1524 2675 1539
rect 175 1477 2675 1492
rect 175 1457 200 1477
rect 220 1457 240 1477
rect 260 1457 280 1477
rect 300 1457 320 1477
rect 340 1457 360 1477
rect 380 1457 400 1477
rect 420 1457 440 1477
rect 460 1457 480 1477
rect 500 1457 520 1477
rect 540 1457 560 1477
rect 580 1457 600 1477
rect 620 1457 640 1477
rect 660 1457 680 1477
rect 700 1457 720 1477
rect 740 1457 760 1477
rect 780 1457 800 1477
rect 820 1457 840 1477
rect 860 1457 880 1477
rect 900 1457 920 1477
rect 940 1457 960 1477
rect 980 1457 1000 1477
rect 1020 1457 1040 1477
rect 1060 1457 1080 1477
rect 1100 1457 1120 1477
rect 1140 1457 1160 1477
rect 1180 1457 1200 1477
rect 1220 1457 1240 1477
rect 1260 1457 1280 1477
rect 1300 1457 1320 1477
rect 1340 1457 1360 1477
rect 1380 1457 1400 1477
rect 1420 1457 1440 1477
rect 1460 1457 1480 1477
rect 1500 1457 1520 1477
rect 1540 1457 1560 1477
rect 1580 1457 1600 1477
rect 1620 1457 1640 1477
rect 1660 1457 1680 1477
rect 1700 1457 1720 1477
rect 1740 1457 1760 1477
rect 1780 1457 1800 1477
rect 1820 1457 1840 1477
rect 1860 1457 1880 1477
rect 1900 1457 1920 1477
rect 1940 1457 1960 1477
rect 1980 1457 2000 1477
rect 2020 1457 2040 1477
rect 2060 1457 2080 1477
rect 2100 1457 2120 1477
rect 2140 1457 2160 1477
rect 2180 1457 2200 1477
rect 2220 1457 2240 1477
rect 2260 1457 2280 1477
rect 2300 1457 2320 1477
rect 2340 1457 2360 1477
rect 2380 1457 2400 1477
rect 2420 1457 2440 1477
rect 2460 1457 2480 1477
rect 2500 1457 2520 1477
rect 2540 1457 2560 1477
rect 2580 1457 2600 1477
rect 2620 1457 2640 1477
rect 2660 1457 2675 1477
rect 175 1442 2675 1457
rect 175 1395 2675 1410
rect 175 1375 200 1395
rect 220 1375 240 1395
rect 260 1375 280 1395
rect 300 1375 320 1395
rect 340 1375 360 1395
rect 380 1375 400 1395
rect 420 1375 440 1395
rect 460 1375 480 1395
rect 500 1375 520 1395
rect 540 1375 560 1395
rect 580 1375 600 1395
rect 620 1375 640 1395
rect 660 1375 680 1395
rect 700 1375 720 1395
rect 740 1375 760 1395
rect 780 1375 800 1395
rect 820 1375 840 1395
rect 860 1375 880 1395
rect 900 1375 920 1395
rect 940 1375 960 1395
rect 980 1375 1000 1395
rect 1020 1375 1040 1395
rect 1060 1375 1080 1395
rect 1100 1375 1120 1395
rect 1140 1375 1160 1395
rect 1180 1375 1200 1395
rect 1220 1375 1240 1395
rect 1260 1375 1280 1395
rect 1300 1375 1320 1395
rect 1340 1375 1360 1395
rect 1380 1375 1400 1395
rect 1420 1375 1440 1395
rect 1460 1375 1480 1395
rect 1500 1375 1520 1395
rect 1540 1375 1560 1395
rect 1580 1375 1600 1395
rect 1620 1375 1640 1395
rect 1660 1375 1680 1395
rect 1700 1375 1720 1395
rect 1740 1375 1760 1395
rect 1780 1375 1800 1395
rect 1820 1375 1840 1395
rect 1860 1375 1880 1395
rect 1900 1375 1920 1395
rect 1940 1375 1960 1395
rect 1980 1375 2000 1395
rect 2020 1375 2040 1395
rect 2060 1375 2080 1395
rect 2100 1375 2120 1395
rect 2140 1375 2160 1395
rect 2180 1375 2200 1395
rect 2220 1375 2240 1395
rect 2260 1375 2280 1395
rect 2300 1375 2320 1395
rect 2340 1375 2360 1395
rect 2380 1375 2400 1395
rect 2420 1375 2440 1395
rect 2460 1375 2480 1395
rect 2500 1375 2520 1395
rect 2540 1375 2560 1395
rect 2580 1375 2600 1395
rect 2620 1375 2640 1395
rect 2660 1375 2675 1395
rect 175 1360 2675 1375
rect 175 1313 2675 1328
rect 175 1293 200 1313
rect 220 1293 240 1313
rect 260 1293 280 1313
rect 300 1293 320 1313
rect 340 1293 360 1313
rect 380 1293 400 1313
rect 420 1293 440 1313
rect 460 1293 480 1313
rect 500 1293 520 1313
rect 540 1293 560 1313
rect 580 1293 600 1313
rect 620 1293 640 1313
rect 660 1293 680 1313
rect 700 1293 720 1313
rect 740 1293 760 1313
rect 780 1293 800 1313
rect 820 1293 840 1313
rect 860 1293 880 1313
rect 900 1293 920 1313
rect 940 1293 960 1313
rect 980 1293 1000 1313
rect 1020 1293 1040 1313
rect 1060 1293 1080 1313
rect 1100 1293 1120 1313
rect 1140 1293 1160 1313
rect 1180 1293 1200 1313
rect 1220 1293 1240 1313
rect 1260 1293 1280 1313
rect 1300 1293 1320 1313
rect 1340 1293 1360 1313
rect 1380 1293 1400 1313
rect 1420 1293 1440 1313
rect 1460 1293 1480 1313
rect 1500 1293 1520 1313
rect 1540 1293 1560 1313
rect 1580 1293 1600 1313
rect 1620 1293 1640 1313
rect 1660 1293 1680 1313
rect 1700 1293 1720 1313
rect 1740 1293 1760 1313
rect 1780 1293 1800 1313
rect 1820 1293 1840 1313
rect 1860 1293 1880 1313
rect 1900 1293 1920 1313
rect 1940 1293 1960 1313
rect 1980 1293 2000 1313
rect 2020 1293 2040 1313
rect 2060 1293 2080 1313
rect 2100 1293 2120 1313
rect 2140 1293 2160 1313
rect 2180 1293 2200 1313
rect 2220 1293 2240 1313
rect 2260 1293 2280 1313
rect 2300 1293 2320 1313
rect 2340 1293 2360 1313
rect 2380 1293 2400 1313
rect 2420 1293 2440 1313
rect 2460 1293 2480 1313
rect 2500 1293 2520 1313
rect 2540 1293 2560 1313
rect 2580 1293 2600 1313
rect 2620 1293 2640 1313
rect 2660 1293 2675 1313
rect 175 1278 2675 1293
rect 175 1231 2675 1246
rect 175 1211 200 1231
rect 220 1211 240 1231
rect 260 1211 280 1231
rect 300 1211 320 1231
rect 340 1211 360 1231
rect 380 1211 400 1231
rect 420 1211 440 1231
rect 460 1211 480 1231
rect 500 1211 520 1231
rect 540 1211 560 1231
rect 580 1211 600 1231
rect 620 1211 640 1231
rect 660 1211 680 1231
rect 700 1211 720 1231
rect 740 1211 760 1231
rect 780 1211 800 1231
rect 820 1211 840 1231
rect 860 1211 880 1231
rect 900 1211 920 1231
rect 940 1211 960 1231
rect 980 1211 1000 1231
rect 1020 1211 1040 1231
rect 1060 1211 1080 1231
rect 1100 1211 1120 1231
rect 1140 1211 1160 1231
rect 1180 1211 1200 1231
rect 1220 1211 1240 1231
rect 1260 1211 1280 1231
rect 1300 1211 1320 1231
rect 1340 1211 1360 1231
rect 1380 1211 1400 1231
rect 1420 1211 1440 1231
rect 1460 1211 1480 1231
rect 1500 1211 1520 1231
rect 1540 1211 1560 1231
rect 1580 1211 1600 1231
rect 1620 1211 1640 1231
rect 1660 1211 1680 1231
rect 1700 1211 1720 1231
rect 1740 1211 1760 1231
rect 1780 1211 1800 1231
rect 1820 1211 1840 1231
rect 1860 1211 1880 1231
rect 1900 1211 1920 1231
rect 1940 1211 1960 1231
rect 1980 1211 2000 1231
rect 2020 1211 2040 1231
rect 2060 1211 2080 1231
rect 2100 1211 2120 1231
rect 2140 1211 2160 1231
rect 2180 1211 2200 1231
rect 2220 1211 2240 1231
rect 2260 1211 2280 1231
rect 2300 1211 2320 1231
rect 2340 1211 2360 1231
rect 2380 1211 2400 1231
rect 2420 1211 2440 1231
rect 2460 1211 2480 1231
rect 2500 1211 2520 1231
rect 2540 1211 2560 1231
rect 2580 1211 2600 1231
rect 2620 1211 2640 1231
rect 2660 1211 2675 1231
rect 175 1196 2675 1211
rect 175 1149 2675 1164
rect 175 1129 200 1149
rect 220 1129 240 1149
rect 260 1129 280 1149
rect 300 1129 320 1149
rect 340 1129 360 1149
rect 380 1129 400 1149
rect 420 1129 440 1149
rect 460 1129 480 1149
rect 500 1129 520 1149
rect 540 1129 560 1149
rect 580 1129 600 1149
rect 620 1129 640 1149
rect 660 1129 680 1149
rect 700 1129 720 1149
rect 740 1129 760 1149
rect 780 1129 800 1149
rect 820 1129 840 1149
rect 860 1129 880 1149
rect 900 1129 920 1149
rect 940 1129 960 1149
rect 980 1129 1000 1149
rect 1020 1129 1040 1149
rect 1060 1129 1080 1149
rect 1100 1129 1120 1149
rect 1140 1129 1160 1149
rect 1180 1129 1200 1149
rect 1220 1129 1240 1149
rect 1260 1129 1280 1149
rect 1300 1129 1320 1149
rect 1340 1129 1360 1149
rect 1380 1129 1400 1149
rect 1420 1129 1440 1149
rect 1460 1129 1480 1149
rect 1500 1129 1520 1149
rect 1540 1129 1560 1149
rect 1580 1129 1600 1149
rect 1620 1129 1640 1149
rect 1660 1129 1680 1149
rect 1700 1129 1720 1149
rect 1740 1129 1760 1149
rect 1780 1129 1800 1149
rect 1820 1129 1840 1149
rect 1860 1129 1880 1149
rect 1900 1129 1920 1149
rect 1940 1129 1960 1149
rect 1980 1129 2000 1149
rect 2020 1129 2040 1149
rect 2060 1129 2080 1149
rect 2100 1129 2120 1149
rect 2140 1129 2160 1149
rect 2180 1129 2200 1149
rect 2220 1129 2240 1149
rect 2260 1129 2280 1149
rect 2300 1129 2320 1149
rect 2340 1129 2360 1149
rect 2380 1129 2400 1149
rect 2420 1129 2440 1149
rect 2460 1129 2480 1149
rect 2500 1129 2520 1149
rect 2540 1129 2560 1149
rect 2580 1129 2600 1149
rect 2620 1129 2640 1149
rect 2660 1129 2675 1149
rect 175 1114 2675 1129
rect 175 1067 2675 1082
rect 175 1047 200 1067
rect 220 1047 240 1067
rect 260 1047 280 1067
rect 300 1047 320 1067
rect 340 1047 360 1067
rect 380 1047 400 1067
rect 420 1047 440 1067
rect 460 1047 480 1067
rect 500 1047 520 1067
rect 540 1047 560 1067
rect 580 1047 600 1067
rect 620 1047 640 1067
rect 660 1047 680 1067
rect 700 1047 720 1067
rect 740 1047 760 1067
rect 780 1047 800 1067
rect 820 1047 840 1067
rect 860 1047 880 1067
rect 900 1047 920 1067
rect 940 1047 960 1067
rect 980 1047 1000 1067
rect 1020 1047 1040 1067
rect 1060 1047 1080 1067
rect 1100 1047 1120 1067
rect 1140 1047 1160 1067
rect 1180 1047 1200 1067
rect 1220 1047 1240 1067
rect 1260 1047 1280 1067
rect 1300 1047 1320 1067
rect 1340 1047 1360 1067
rect 1380 1047 1400 1067
rect 1420 1047 1440 1067
rect 1460 1047 1480 1067
rect 1500 1047 1520 1067
rect 1540 1047 1560 1067
rect 1580 1047 1600 1067
rect 1620 1047 1640 1067
rect 1660 1047 1680 1067
rect 1700 1047 1720 1067
rect 1740 1047 1760 1067
rect 1780 1047 1800 1067
rect 1820 1047 1840 1067
rect 1860 1047 1880 1067
rect 1900 1047 1920 1067
rect 1940 1047 1960 1067
rect 1980 1047 2000 1067
rect 2020 1047 2040 1067
rect 2060 1047 2080 1067
rect 2100 1047 2120 1067
rect 2140 1047 2160 1067
rect 2180 1047 2200 1067
rect 2220 1047 2240 1067
rect 2260 1047 2280 1067
rect 2300 1047 2320 1067
rect 2340 1047 2360 1067
rect 2380 1047 2400 1067
rect 2420 1047 2440 1067
rect 2460 1047 2480 1067
rect 2500 1047 2520 1067
rect 2540 1047 2560 1067
rect 2580 1047 2600 1067
rect 2620 1047 2640 1067
rect 2660 1047 2675 1067
rect 175 1032 2675 1047
rect 175 985 2675 1000
rect 175 965 200 985
rect 220 965 240 985
rect 260 965 280 985
rect 300 965 320 985
rect 340 965 360 985
rect 380 965 400 985
rect 420 965 440 985
rect 460 965 480 985
rect 500 965 520 985
rect 540 965 560 985
rect 580 965 600 985
rect 620 965 640 985
rect 660 965 680 985
rect 700 965 720 985
rect 740 965 760 985
rect 780 965 800 985
rect 820 965 840 985
rect 860 965 880 985
rect 900 965 920 985
rect 940 965 960 985
rect 980 965 1000 985
rect 1020 965 1040 985
rect 1060 965 1080 985
rect 1100 965 1120 985
rect 1140 965 1160 985
rect 1180 965 1200 985
rect 1220 965 1240 985
rect 1260 965 1280 985
rect 1300 965 1320 985
rect 1340 965 1360 985
rect 1380 965 1400 985
rect 1420 965 1440 985
rect 1460 965 1480 985
rect 1500 965 1520 985
rect 1540 965 1560 985
rect 1580 965 1600 985
rect 1620 965 1640 985
rect 1660 965 1680 985
rect 1700 965 1720 985
rect 1740 965 1760 985
rect 1780 965 1800 985
rect 1820 965 1840 985
rect 1860 965 1880 985
rect 1900 965 1920 985
rect 1940 965 1960 985
rect 1980 965 2000 985
rect 2020 965 2040 985
rect 2060 965 2080 985
rect 2100 965 2120 985
rect 2140 965 2160 985
rect 2180 965 2200 985
rect 2220 965 2240 985
rect 2260 965 2280 985
rect 2300 965 2320 985
rect 2340 965 2360 985
rect 2380 965 2400 985
rect 2420 965 2440 985
rect 2460 965 2480 985
rect 2500 965 2520 985
rect 2540 965 2560 985
rect 2580 965 2600 985
rect 2620 965 2640 985
rect 2660 965 2675 985
rect 175 950 2675 965
rect 175 903 2675 918
rect 175 883 200 903
rect 220 883 240 903
rect 260 883 280 903
rect 300 883 320 903
rect 340 883 360 903
rect 380 883 400 903
rect 420 883 440 903
rect 460 883 480 903
rect 500 883 520 903
rect 540 883 560 903
rect 580 883 600 903
rect 620 883 640 903
rect 660 883 680 903
rect 700 883 720 903
rect 740 883 760 903
rect 780 883 800 903
rect 820 883 840 903
rect 860 883 880 903
rect 900 883 920 903
rect 940 883 960 903
rect 980 883 1000 903
rect 1020 883 1040 903
rect 1060 883 1080 903
rect 1100 883 1120 903
rect 1140 883 1160 903
rect 1180 883 1200 903
rect 1220 883 1240 903
rect 1260 883 1280 903
rect 1300 883 1320 903
rect 1340 883 1360 903
rect 1380 883 1400 903
rect 1420 883 1440 903
rect 1460 883 1480 903
rect 1500 883 1520 903
rect 1540 883 1560 903
rect 1580 883 1600 903
rect 1620 883 1640 903
rect 1660 883 1680 903
rect 1700 883 1720 903
rect 1740 883 1760 903
rect 1780 883 1800 903
rect 1820 883 1840 903
rect 1860 883 1880 903
rect 1900 883 1920 903
rect 1940 883 1960 903
rect 1980 883 2000 903
rect 2020 883 2040 903
rect 2060 883 2080 903
rect 2100 883 2120 903
rect 2140 883 2160 903
rect 2180 883 2200 903
rect 2220 883 2240 903
rect 2260 883 2280 903
rect 2300 883 2320 903
rect 2340 883 2360 903
rect 2380 883 2400 903
rect 2420 883 2440 903
rect 2460 883 2480 903
rect 2500 883 2520 903
rect 2540 883 2560 903
rect 2580 883 2600 903
rect 2620 883 2640 903
rect 2660 883 2675 903
rect 175 868 2675 883
rect 175 821 2675 836
rect 175 801 200 821
rect 220 801 240 821
rect 260 801 280 821
rect 300 801 320 821
rect 340 801 360 821
rect 380 801 400 821
rect 420 801 440 821
rect 460 801 480 821
rect 500 801 520 821
rect 540 801 560 821
rect 580 801 600 821
rect 620 801 640 821
rect 660 801 680 821
rect 700 801 720 821
rect 740 801 760 821
rect 780 801 800 821
rect 820 801 840 821
rect 860 801 880 821
rect 900 801 920 821
rect 940 801 960 821
rect 980 801 1000 821
rect 1020 801 1040 821
rect 1060 801 1080 821
rect 1100 801 1120 821
rect 1140 801 1160 821
rect 1180 801 1200 821
rect 1220 801 1240 821
rect 1260 801 1280 821
rect 1300 801 1320 821
rect 1340 801 1360 821
rect 1380 801 1400 821
rect 1420 801 1440 821
rect 1460 801 1480 821
rect 1500 801 1520 821
rect 1540 801 1560 821
rect 1580 801 1600 821
rect 1620 801 1640 821
rect 1660 801 1680 821
rect 1700 801 1720 821
rect 1740 801 1760 821
rect 1780 801 1800 821
rect 1820 801 1840 821
rect 1860 801 1880 821
rect 1900 801 1920 821
rect 1940 801 1960 821
rect 1980 801 2000 821
rect 2020 801 2040 821
rect 2060 801 2080 821
rect 2100 801 2120 821
rect 2140 801 2160 821
rect 2180 801 2200 821
rect 2220 801 2240 821
rect 2260 801 2280 821
rect 2300 801 2320 821
rect 2340 801 2360 821
rect 2380 801 2400 821
rect 2420 801 2440 821
rect 2460 801 2480 821
rect 2500 801 2520 821
rect 2540 801 2560 821
rect 2580 801 2600 821
rect 2620 801 2640 821
rect 2660 801 2675 821
rect 175 786 2675 801
rect 175 739 2675 754
rect 175 719 200 739
rect 220 719 240 739
rect 260 719 280 739
rect 300 719 320 739
rect 340 719 360 739
rect 380 719 400 739
rect 420 719 440 739
rect 460 719 480 739
rect 500 719 520 739
rect 540 719 560 739
rect 580 719 600 739
rect 620 719 640 739
rect 660 719 680 739
rect 700 719 720 739
rect 740 719 760 739
rect 780 719 800 739
rect 820 719 840 739
rect 860 719 880 739
rect 900 719 920 739
rect 940 719 960 739
rect 980 719 1000 739
rect 1020 719 1040 739
rect 1060 719 1080 739
rect 1100 719 1120 739
rect 1140 719 1160 739
rect 1180 719 1200 739
rect 1220 719 1240 739
rect 1260 719 1280 739
rect 1300 719 1320 739
rect 1340 719 1360 739
rect 1380 719 1400 739
rect 1420 719 1440 739
rect 1460 719 1480 739
rect 1500 719 1520 739
rect 1540 719 1560 739
rect 1580 719 1600 739
rect 1620 719 1640 739
rect 1660 719 1680 739
rect 1700 719 1720 739
rect 1740 719 1760 739
rect 1780 719 1800 739
rect 1820 719 1840 739
rect 1860 719 1880 739
rect 1900 719 1920 739
rect 1940 719 1960 739
rect 1980 719 2000 739
rect 2020 719 2040 739
rect 2060 719 2080 739
rect 2100 719 2120 739
rect 2140 719 2160 739
rect 2180 719 2200 739
rect 2220 719 2240 739
rect 2260 719 2280 739
rect 2300 719 2320 739
rect 2340 719 2360 739
rect 2380 719 2400 739
rect 2420 719 2440 739
rect 2460 719 2480 739
rect 2500 719 2520 739
rect 2540 719 2560 739
rect 2580 719 2600 739
rect 2620 719 2640 739
rect 2660 719 2675 739
rect 175 704 2675 719
rect 175 657 2675 672
rect 175 637 200 657
rect 220 637 240 657
rect 260 637 280 657
rect 300 637 320 657
rect 340 637 360 657
rect 380 637 400 657
rect 420 637 440 657
rect 460 637 480 657
rect 500 637 520 657
rect 540 637 560 657
rect 580 637 600 657
rect 620 637 640 657
rect 660 637 680 657
rect 700 637 720 657
rect 740 637 760 657
rect 780 637 800 657
rect 820 637 840 657
rect 860 637 880 657
rect 900 637 920 657
rect 940 637 960 657
rect 980 637 1000 657
rect 1020 637 1040 657
rect 1060 637 1080 657
rect 1100 637 1120 657
rect 1140 637 1160 657
rect 1180 637 1200 657
rect 1220 637 1240 657
rect 1260 637 1280 657
rect 1300 637 1320 657
rect 1340 637 1360 657
rect 1380 637 1400 657
rect 1420 637 1440 657
rect 1460 637 1480 657
rect 1500 637 1520 657
rect 1540 637 1560 657
rect 1580 637 1600 657
rect 1620 637 1640 657
rect 1660 637 1680 657
rect 1700 637 1720 657
rect 1740 637 1760 657
rect 1780 637 1800 657
rect 1820 637 1840 657
rect 1860 637 1880 657
rect 1900 637 1920 657
rect 1940 637 1960 657
rect 1980 637 2000 657
rect 2020 637 2040 657
rect 2060 637 2080 657
rect 2100 637 2120 657
rect 2140 637 2160 657
rect 2180 637 2200 657
rect 2220 637 2240 657
rect 2260 637 2280 657
rect 2300 637 2320 657
rect 2340 637 2360 657
rect 2380 637 2400 657
rect 2420 637 2440 657
rect 2460 637 2480 657
rect 2500 637 2520 657
rect 2540 637 2560 657
rect 2580 637 2600 657
rect 2620 637 2640 657
rect 2660 637 2675 657
rect 175 622 2675 637
rect 175 575 2675 590
rect 175 555 200 575
rect 220 555 240 575
rect 260 555 280 575
rect 300 555 320 575
rect 340 555 360 575
rect 380 555 400 575
rect 420 555 440 575
rect 460 555 480 575
rect 500 555 520 575
rect 540 555 560 575
rect 580 555 600 575
rect 620 555 640 575
rect 660 555 680 575
rect 700 555 720 575
rect 740 555 760 575
rect 780 555 800 575
rect 820 555 840 575
rect 860 555 880 575
rect 900 555 920 575
rect 940 555 960 575
rect 980 555 1000 575
rect 1020 555 1040 575
rect 1060 555 1080 575
rect 1100 555 1120 575
rect 1140 555 1160 575
rect 1180 555 1200 575
rect 1220 555 1240 575
rect 1260 555 1280 575
rect 1300 555 1320 575
rect 1340 555 1360 575
rect 1380 555 1400 575
rect 1420 555 1440 575
rect 1460 555 1480 575
rect 1500 555 1520 575
rect 1540 555 1560 575
rect 1580 555 1600 575
rect 1620 555 1640 575
rect 1660 555 1680 575
rect 1700 555 1720 575
rect 1740 555 1760 575
rect 1780 555 1800 575
rect 1820 555 1840 575
rect 1860 555 1880 575
rect 1900 555 1920 575
rect 1940 555 1960 575
rect 1980 555 2000 575
rect 2020 555 2040 575
rect 2060 555 2080 575
rect 2100 555 2120 575
rect 2140 555 2160 575
rect 2180 555 2200 575
rect 2220 555 2240 575
rect 2260 555 2280 575
rect 2300 555 2320 575
rect 2340 555 2360 575
rect 2380 555 2400 575
rect 2420 555 2440 575
rect 2460 555 2480 575
rect 2500 555 2520 575
rect 2540 555 2560 575
rect 2580 555 2600 575
rect 2620 555 2640 575
rect 2660 555 2675 575
rect 175 540 2675 555
rect 175 493 2675 508
rect 175 473 200 493
rect 220 473 240 493
rect 260 473 280 493
rect 300 473 320 493
rect 340 473 360 493
rect 380 473 400 493
rect 420 473 440 493
rect 460 473 480 493
rect 500 473 520 493
rect 540 473 560 493
rect 580 473 600 493
rect 620 473 640 493
rect 660 473 680 493
rect 700 473 720 493
rect 740 473 760 493
rect 780 473 800 493
rect 820 473 840 493
rect 860 473 880 493
rect 900 473 920 493
rect 940 473 960 493
rect 980 473 1000 493
rect 1020 473 1040 493
rect 1060 473 1080 493
rect 1100 473 1120 493
rect 1140 473 1160 493
rect 1180 473 1200 493
rect 1220 473 1240 493
rect 1260 473 1280 493
rect 1300 473 1320 493
rect 1340 473 1360 493
rect 1380 473 1400 493
rect 1420 473 1440 493
rect 1460 473 1480 493
rect 1500 473 1520 493
rect 1540 473 1560 493
rect 1580 473 1600 493
rect 1620 473 1640 493
rect 1660 473 1680 493
rect 1700 473 1720 493
rect 1740 473 1760 493
rect 1780 473 1800 493
rect 1820 473 1840 493
rect 1860 473 1880 493
rect 1900 473 1920 493
rect 1940 473 1960 493
rect 1980 473 2000 493
rect 2020 473 2040 493
rect 2060 473 2080 493
rect 2100 473 2120 493
rect 2140 473 2160 493
rect 2180 473 2200 493
rect 2220 473 2240 493
rect 2260 473 2280 493
rect 2300 473 2320 493
rect 2340 473 2360 493
rect 2380 473 2400 493
rect 2420 473 2440 493
rect 2460 473 2480 493
rect 2500 473 2520 493
rect 2540 473 2560 493
rect 2580 473 2600 493
rect 2620 473 2640 493
rect 2660 473 2675 493
rect 175 458 2675 473
rect 175 411 2675 426
rect 175 391 200 411
rect 220 391 240 411
rect 260 391 280 411
rect 300 391 320 411
rect 340 391 360 411
rect 380 391 400 411
rect 420 391 440 411
rect 460 391 480 411
rect 500 391 520 411
rect 540 391 560 411
rect 580 391 600 411
rect 620 391 640 411
rect 660 391 680 411
rect 700 391 720 411
rect 740 391 760 411
rect 780 391 800 411
rect 820 391 840 411
rect 860 391 880 411
rect 900 391 920 411
rect 940 391 960 411
rect 980 391 1000 411
rect 1020 391 1040 411
rect 1060 391 1080 411
rect 1100 391 1120 411
rect 1140 391 1160 411
rect 1180 391 1200 411
rect 1220 391 1240 411
rect 1260 391 1280 411
rect 1300 391 1320 411
rect 1340 391 1360 411
rect 1380 391 1400 411
rect 1420 391 1440 411
rect 1460 391 1480 411
rect 1500 391 1520 411
rect 1540 391 1560 411
rect 1580 391 1600 411
rect 1620 391 1640 411
rect 1660 391 1680 411
rect 1700 391 1720 411
rect 1740 391 1760 411
rect 1780 391 1800 411
rect 1820 391 1840 411
rect 1860 391 1880 411
rect 1900 391 1920 411
rect 1940 391 1960 411
rect 1980 391 2000 411
rect 2020 391 2040 411
rect 2060 391 2080 411
rect 2100 391 2120 411
rect 2140 391 2160 411
rect 2180 391 2200 411
rect 2220 391 2240 411
rect 2260 391 2280 411
rect 2300 391 2320 411
rect 2340 391 2360 411
rect 2380 391 2400 411
rect 2420 391 2440 411
rect 2460 391 2480 411
rect 2500 391 2520 411
rect 2540 391 2560 411
rect 2580 391 2600 411
rect 2620 391 2640 411
rect 2660 391 2675 411
rect 175 376 2675 391
rect 175 329 2675 344
rect 175 309 200 329
rect 220 309 240 329
rect 260 309 280 329
rect 300 309 320 329
rect 340 309 360 329
rect 380 309 400 329
rect 420 309 440 329
rect 460 309 480 329
rect 500 309 520 329
rect 540 309 560 329
rect 580 309 600 329
rect 620 309 640 329
rect 660 309 680 329
rect 700 309 720 329
rect 740 309 760 329
rect 780 309 800 329
rect 820 309 840 329
rect 860 309 880 329
rect 900 309 920 329
rect 940 309 960 329
rect 980 309 1000 329
rect 1020 309 1040 329
rect 1060 309 1080 329
rect 1100 309 1120 329
rect 1140 309 1160 329
rect 1180 309 1200 329
rect 1220 309 1240 329
rect 1260 309 1280 329
rect 1300 309 1320 329
rect 1340 309 1360 329
rect 1380 309 1400 329
rect 1420 309 1440 329
rect 1460 309 1480 329
rect 1500 309 1520 329
rect 1540 309 1560 329
rect 1580 309 1600 329
rect 1620 309 1640 329
rect 1660 309 1680 329
rect 1700 309 1720 329
rect 1740 309 1760 329
rect 1780 309 1800 329
rect 1820 309 1840 329
rect 1860 309 1880 329
rect 1900 309 1920 329
rect 1940 309 1960 329
rect 1980 309 2000 329
rect 2020 309 2040 329
rect 2060 309 2080 329
rect 2100 309 2120 329
rect 2140 309 2160 329
rect 2180 309 2200 329
rect 2220 309 2240 329
rect 2260 309 2280 329
rect 2300 309 2320 329
rect 2340 309 2360 329
rect 2380 309 2400 329
rect 2420 309 2440 329
rect 2460 309 2480 329
rect 2500 309 2520 329
rect 2540 309 2560 329
rect 2580 309 2600 329
rect 2620 309 2640 329
rect 2660 309 2675 329
rect 175 294 2675 309
rect 175 247 2675 262
rect 175 227 200 247
rect 220 227 240 247
rect 260 227 280 247
rect 300 227 320 247
rect 340 227 360 247
rect 380 227 400 247
rect 420 227 440 247
rect 460 227 480 247
rect 500 227 520 247
rect 540 227 560 247
rect 580 227 600 247
rect 620 227 640 247
rect 660 227 680 247
rect 700 227 720 247
rect 740 227 760 247
rect 780 227 800 247
rect 820 227 840 247
rect 860 227 880 247
rect 900 227 920 247
rect 940 227 960 247
rect 980 227 1000 247
rect 1020 227 1040 247
rect 1060 227 1080 247
rect 1100 227 1120 247
rect 1140 227 1160 247
rect 1180 227 1200 247
rect 1220 227 1240 247
rect 1260 227 1280 247
rect 1300 227 1320 247
rect 1340 227 1360 247
rect 1380 227 1400 247
rect 1420 227 1440 247
rect 1460 227 1480 247
rect 1500 227 1520 247
rect 1540 227 1560 247
rect 1580 227 1600 247
rect 1620 227 1640 247
rect 1660 227 1680 247
rect 1700 227 1720 247
rect 1740 227 1760 247
rect 1780 227 1800 247
rect 1820 227 1840 247
rect 1860 227 1880 247
rect 1900 227 1920 247
rect 1940 227 1960 247
rect 1980 227 2000 247
rect 2020 227 2040 247
rect 2060 227 2080 247
rect 2100 227 2120 247
rect 2140 227 2160 247
rect 2180 227 2200 247
rect 2220 227 2240 247
rect 2260 227 2280 247
rect 2300 227 2320 247
rect 2340 227 2360 247
rect 2380 227 2400 247
rect 2420 227 2440 247
rect 2460 227 2480 247
rect 2500 227 2520 247
rect 2540 227 2560 247
rect 2580 227 2600 247
rect 2620 227 2640 247
rect 2660 227 2675 247
rect 175 212 2675 227
rect 175 165 2675 180
rect 175 145 200 165
rect 220 145 240 165
rect 260 145 280 165
rect 300 145 320 165
rect 340 145 360 165
rect 380 145 400 165
rect 420 145 440 165
rect 460 145 480 165
rect 500 145 520 165
rect 540 145 560 165
rect 580 145 600 165
rect 620 145 640 165
rect 660 145 680 165
rect 700 145 720 165
rect 740 145 760 165
rect 780 145 800 165
rect 820 145 840 165
rect 860 145 880 165
rect 900 145 920 165
rect 940 145 960 165
rect 980 145 1000 165
rect 1020 145 1040 165
rect 1060 145 1080 165
rect 1100 145 1120 165
rect 1140 145 1160 165
rect 1180 145 1200 165
rect 1220 145 1240 165
rect 1260 145 1280 165
rect 1300 145 1320 165
rect 1340 145 1360 165
rect 1380 145 1400 165
rect 1420 145 1440 165
rect 1460 145 1480 165
rect 1500 145 1520 165
rect 1540 145 1560 165
rect 1580 145 1600 165
rect 1620 145 1640 165
rect 1660 145 1680 165
rect 1700 145 1720 165
rect 1740 145 1760 165
rect 1780 145 1800 165
rect 1820 145 1840 165
rect 1860 145 1880 165
rect 1900 145 1920 165
rect 1940 145 1960 165
rect 1980 145 2000 165
rect 2020 145 2040 165
rect 2060 145 2080 165
rect 2100 145 2120 165
rect 2140 145 2160 165
rect 2180 145 2200 165
rect 2220 145 2240 165
rect 2260 145 2280 165
rect 2300 145 2320 165
rect 2340 145 2360 165
rect 2380 145 2400 165
rect 2420 145 2440 165
rect 2460 145 2480 165
rect 2500 145 2520 165
rect 2540 145 2560 165
rect 2580 145 2600 165
rect 2620 145 2640 165
rect 2660 145 2675 165
rect 175 135 2675 145
rect 105 -50 2605 -40
rect 105 -70 120 -50
rect 140 -70 160 -50
rect 180 -70 200 -50
rect 220 -70 240 -50
rect 260 -70 280 -50
rect 300 -70 320 -50
rect 340 -70 360 -50
rect 380 -70 400 -50
rect 420 -70 440 -50
rect 460 -70 480 -50
rect 500 -70 520 -50
rect 540 -70 560 -50
rect 580 -70 600 -50
rect 620 -70 640 -50
rect 660 -70 680 -50
rect 700 -70 720 -50
rect 740 -70 760 -50
rect 780 -70 800 -50
rect 820 -70 840 -50
rect 860 -70 880 -50
rect 900 -70 920 -50
rect 940 -70 960 -50
rect 980 -70 1000 -50
rect 1020 -70 1040 -50
rect 1060 -70 1080 -50
rect 1100 -70 1120 -50
rect 1140 -70 1160 -50
rect 1180 -70 1200 -50
rect 1220 -70 1240 -50
rect 1260 -70 1280 -50
rect 1300 -70 1320 -50
rect 1340 -70 1360 -50
rect 1380 -70 1400 -50
rect 1420 -70 1440 -50
rect 1460 -70 1480 -50
rect 1500 -70 1520 -50
rect 1540 -70 1560 -50
rect 1580 -70 1600 -50
rect 1620 -70 1640 -50
rect 1660 -70 1680 -50
rect 1700 -70 1720 -50
rect 1740 -70 1760 -50
rect 1780 -70 1800 -50
rect 1820 -70 1840 -50
rect 1860 -70 1880 -50
rect 1900 -70 1920 -50
rect 1940 -70 1960 -50
rect 1980 -70 2000 -50
rect 2020 -70 2040 -50
rect 2060 -70 2080 -50
rect 2100 -70 2120 -50
rect 2140 -70 2160 -50
rect 2180 -70 2200 -50
rect 2220 -70 2240 -50
rect 2260 -70 2280 -50
rect 2300 -70 2320 -50
rect 2340 -70 2360 -50
rect 2380 -70 2400 -50
rect 2420 -70 2440 -50
rect 2460 -70 2480 -50
rect 2500 -70 2520 -50
rect 2540 -70 2560 -50
rect 2590 -70 2605 -50
rect 105 -85 2605 -70
rect 105 -145 2605 -130
rect 105 -165 120 -145
rect 140 -165 160 -145
rect 180 -165 200 -145
rect 220 -165 240 -145
rect 260 -165 280 -145
rect 300 -165 320 -145
rect 340 -165 360 -145
rect 380 -165 400 -145
rect 420 -165 440 -145
rect 460 -165 480 -145
rect 500 -165 520 -145
rect 540 -165 560 -145
rect 580 -165 600 -145
rect 620 -165 640 -145
rect 660 -165 680 -145
rect 700 -165 720 -145
rect 740 -165 760 -145
rect 780 -165 800 -145
rect 820 -165 840 -145
rect 860 -165 880 -145
rect 900 -165 920 -145
rect 940 -165 960 -145
rect 980 -165 1000 -145
rect 1020 -165 1040 -145
rect 1060 -165 1080 -145
rect 1100 -165 1120 -145
rect 1140 -165 1160 -145
rect 1180 -165 1200 -145
rect 1220 -165 1240 -145
rect 1260 -165 1280 -145
rect 1300 -165 1320 -145
rect 1340 -165 1360 -145
rect 1380 -165 1400 -145
rect 1420 -165 1440 -145
rect 1460 -165 1480 -145
rect 1500 -165 1520 -145
rect 1540 -165 1560 -145
rect 1580 -165 1600 -145
rect 1620 -165 1640 -145
rect 1660 -165 1680 -145
rect 1700 -165 1720 -145
rect 1740 -165 1760 -145
rect 1780 -165 1800 -145
rect 1820 -165 1840 -145
rect 1860 -165 1880 -145
rect 1900 -165 1920 -145
rect 1940 -165 1960 -145
rect 1980 -165 2000 -145
rect 2020 -165 2040 -145
rect 2060 -165 2080 -145
rect 2100 -165 2120 -145
rect 2140 -165 2160 -145
rect 2180 -165 2200 -145
rect 2220 -165 2240 -145
rect 2260 -165 2280 -145
rect 2300 -165 2320 -145
rect 2340 -165 2360 -145
rect 2380 -165 2400 -145
rect 2420 -165 2440 -145
rect 2460 -165 2480 -145
rect 2500 -165 2520 -145
rect 2540 -165 2560 -145
rect 2590 -165 2605 -145
rect 105 -180 2605 -165
rect 105 -240 2605 -225
rect 105 -260 120 -240
rect 140 -260 160 -240
rect 180 -260 200 -240
rect 220 -260 240 -240
rect 260 -260 280 -240
rect 300 -260 320 -240
rect 340 -260 360 -240
rect 380 -260 400 -240
rect 420 -260 440 -240
rect 460 -260 480 -240
rect 500 -260 520 -240
rect 540 -260 560 -240
rect 580 -260 600 -240
rect 620 -260 640 -240
rect 660 -260 680 -240
rect 700 -260 720 -240
rect 740 -260 760 -240
rect 780 -260 800 -240
rect 820 -260 840 -240
rect 860 -260 880 -240
rect 900 -260 920 -240
rect 940 -260 960 -240
rect 980 -260 1000 -240
rect 1020 -260 1040 -240
rect 1060 -260 1080 -240
rect 1100 -260 1120 -240
rect 1140 -260 1160 -240
rect 1180 -260 1200 -240
rect 1220 -260 1240 -240
rect 1260 -260 1280 -240
rect 1300 -260 1320 -240
rect 1340 -260 1360 -240
rect 1380 -260 1400 -240
rect 1420 -260 1440 -240
rect 1460 -260 1480 -240
rect 1500 -260 1520 -240
rect 1540 -260 1560 -240
rect 1580 -260 1600 -240
rect 1620 -260 1640 -240
rect 1660 -260 1680 -240
rect 1700 -260 1720 -240
rect 1740 -260 1760 -240
rect 1780 -260 1800 -240
rect 1820 -260 1840 -240
rect 1860 -260 1880 -240
rect 1900 -260 1920 -240
rect 1940 -260 1960 -240
rect 1980 -260 2000 -240
rect 2020 -260 2040 -240
rect 2060 -260 2080 -240
rect 2100 -260 2120 -240
rect 2140 -260 2160 -240
rect 2180 -260 2200 -240
rect 2220 -260 2240 -240
rect 2260 -260 2280 -240
rect 2300 -260 2320 -240
rect 2340 -260 2360 -240
rect 2380 -260 2400 -240
rect 2420 -260 2440 -240
rect 2460 -260 2480 -240
rect 2500 -260 2520 -240
rect 2540 -260 2560 -240
rect 2590 -260 2605 -240
rect 105 -275 2605 -260
rect 105 -335 2605 -320
rect 105 -355 120 -335
rect 140 -355 160 -335
rect 180 -355 200 -335
rect 220 -355 240 -335
rect 260 -355 280 -335
rect 300 -355 320 -335
rect 340 -355 360 -335
rect 380 -355 400 -335
rect 420 -355 440 -335
rect 460 -355 480 -335
rect 500 -355 520 -335
rect 540 -355 560 -335
rect 580 -355 600 -335
rect 620 -355 640 -335
rect 660 -355 680 -335
rect 700 -355 720 -335
rect 740 -355 760 -335
rect 780 -355 800 -335
rect 820 -355 840 -335
rect 860 -355 880 -335
rect 900 -355 920 -335
rect 940 -355 960 -335
rect 980 -355 1000 -335
rect 1020 -355 1040 -335
rect 1060 -355 1080 -335
rect 1100 -355 1120 -335
rect 1140 -355 1160 -335
rect 1180 -355 1200 -335
rect 1220 -355 1240 -335
rect 1260 -355 1280 -335
rect 1300 -355 1320 -335
rect 1340 -355 1360 -335
rect 1380 -355 1400 -335
rect 1420 -355 1440 -335
rect 1460 -355 1480 -335
rect 1500 -355 1520 -335
rect 1540 -355 1560 -335
rect 1580 -355 1600 -335
rect 1620 -355 1640 -335
rect 1660 -355 1680 -335
rect 1700 -355 1720 -335
rect 1740 -355 1760 -335
rect 1780 -355 1800 -335
rect 1820 -355 1840 -335
rect 1860 -355 1880 -335
rect 1900 -355 1920 -335
rect 1940 -355 1960 -335
rect 1980 -355 2000 -335
rect 2020 -355 2040 -335
rect 2060 -355 2080 -335
rect 2100 -355 2120 -335
rect 2140 -355 2160 -335
rect 2180 -355 2200 -335
rect 2220 -355 2240 -335
rect 2260 -355 2280 -335
rect 2300 -355 2320 -335
rect 2340 -355 2360 -335
rect 2380 -355 2400 -335
rect 2420 -355 2440 -335
rect 2460 -355 2480 -335
rect 2500 -355 2520 -335
rect 2540 -355 2560 -335
rect 2590 -355 2605 -335
rect 105 -370 2605 -355
rect 105 -430 2605 -415
rect 105 -450 120 -430
rect 140 -450 160 -430
rect 180 -450 200 -430
rect 220 -450 240 -430
rect 260 -450 280 -430
rect 300 -450 320 -430
rect 340 -450 360 -430
rect 380 -450 400 -430
rect 420 -450 440 -430
rect 460 -450 480 -430
rect 500 -450 520 -430
rect 540 -450 560 -430
rect 580 -450 600 -430
rect 620 -450 640 -430
rect 660 -450 680 -430
rect 700 -450 720 -430
rect 740 -450 760 -430
rect 780 -450 800 -430
rect 820 -450 840 -430
rect 860 -450 880 -430
rect 900 -450 920 -430
rect 940 -450 960 -430
rect 980 -450 1000 -430
rect 1020 -450 1040 -430
rect 1060 -450 1080 -430
rect 1100 -450 1120 -430
rect 1140 -450 1160 -430
rect 1180 -450 1200 -430
rect 1220 -450 1240 -430
rect 1260 -450 1280 -430
rect 1300 -450 1320 -430
rect 1340 -450 1360 -430
rect 1380 -450 1400 -430
rect 1420 -450 1440 -430
rect 1460 -450 1480 -430
rect 1500 -450 1520 -430
rect 1540 -450 1560 -430
rect 1580 -450 1600 -430
rect 1620 -450 1640 -430
rect 1660 -450 1680 -430
rect 1700 -450 1720 -430
rect 1740 -450 1760 -430
rect 1780 -450 1800 -430
rect 1820 -450 1840 -430
rect 1860 -450 1880 -430
rect 1900 -450 1920 -430
rect 1940 -450 1960 -430
rect 1980 -450 2000 -430
rect 2020 -450 2040 -430
rect 2060 -450 2080 -430
rect 2100 -450 2120 -430
rect 2140 -450 2160 -430
rect 2180 -450 2200 -430
rect 2220 -450 2240 -430
rect 2260 -450 2280 -430
rect 2300 -450 2320 -430
rect 2340 -450 2360 -430
rect 2380 -450 2400 -430
rect 2420 -450 2440 -430
rect 2460 -450 2480 -430
rect 2500 -450 2520 -430
rect 2540 -450 2560 -430
rect 2590 -450 2605 -430
rect 105 -465 2605 -450
rect 105 -525 2605 -510
rect 105 -545 120 -525
rect 140 -545 160 -525
rect 180 -545 200 -525
rect 220 -545 240 -525
rect 260 -545 280 -525
rect 300 -545 320 -525
rect 340 -545 360 -525
rect 380 -545 400 -525
rect 420 -545 440 -525
rect 460 -545 480 -525
rect 500 -545 520 -525
rect 540 -545 560 -525
rect 580 -545 600 -525
rect 620 -545 640 -525
rect 660 -545 680 -525
rect 700 -545 720 -525
rect 740 -545 760 -525
rect 780 -545 800 -525
rect 820 -545 840 -525
rect 860 -545 880 -525
rect 900 -545 920 -525
rect 940 -545 960 -525
rect 980 -545 1000 -525
rect 1020 -545 1040 -525
rect 1060 -545 1080 -525
rect 1100 -545 1120 -525
rect 1140 -545 1160 -525
rect 1180 -545 1200 -525
rect 1220 -545 1240 -525
rect 1260 -545 1280 -525
rect 1300 -545 1320 -525
rect 1340 -545 1360 -525
rect 1380 -545 1400 -525
rect 1420 -545 1440 -525
rect 1460 -545 1480 -525
rect 1500 -545 1520 -525
rect 1540 -545 1560 -525
rect 1580 -545 1600 -525
rect 1620 -545 1640 -525
rect 1660 -545 1680 -525
rect 1700 -545 1720 -525
rect 1740 -545 1760 -525
rect 1780 -545 1800 -525
rect 1820 -545 1840 -525
rect 1860 -545 1880 -525
rect 1900 -545 1920 -525
rect 1940 -545 1960 -525
rect 1980 -545 2000 -525
rect 2020 -545 2040 -525
rect 2060 -545 2080 -525
rect 2100 -545 2120 -525
rect 2140 -545 2160 -525
rect 2180 -545 2200 -525
rect 2220 -545 2240 -525
rect 2260 -545 2280 -525
rect 2300 -545 2320 -525
rect 2340 -545 2360 -525
rect 2380 -545 2400 -525
rect 2420 -545 2440 -525
rect 2460 -545 2480 -525
rect 2500 -545 2520 -525
rect 2540 -545 2560 -525
rect 2590 -545 2605 -525
rect 105 -560 2605 -545
rect 105 -620 2605 -605
rect 105 -640 120 -620
rect 140 -640 160 -620
rect 180 -640 200 -620
rect 220 -640 240 -620
rect 260 -640 280 -620
rect 300 -640 320 -620
rect 340 -640 360 -620
rect 380 -640 400 -620
rect 420 -640 440 -620
rect 460 -640 480 -620
rect 500 -640 520 -620
rect 540 -640 560 -620
rect 580 -640 600 -620
rect 620 -640 640 -620
rect 660 -640 680 -620
rect 700 -640 720 -620
rect 740 -640 760 -620
rect 780 -640 800 -620
rect 820 -640 840 -620
rect 860 -640 880 -620
rect 900 -640 920 -620
rect 940 -640 960 -620
rect 980 -640 1000 -620
rect 1020 -640 1040 -620
rect 1060 -640 1080 -620
rect 1100 -640 1120 -620
rect 1140 -640 1160 -620
rect 1180 -640 1200 -620
rect 1220 -640 1240 -620
rect 1260 -640 1280 -620
rect 1300 -640 1320 -620
rect 1340 -640 1360 -620
rect 1380 -640 1400 -620
rect 1420 -640 1440 -620
rect 1460 -640 1480 -620
rect 1500 -640 1520 -620
rect 1540 -640 1560 -620
rect 1580 -640 1600 -620
rect 1620 -640 1640 -620
rect 1660 -640 1680 -620
rect 1700 -640 1720 -620
rect 1740 -640 1760 -620
rect 1780 -640 1800 -620
rect 1820 -640 1840 -620
rect 1860 -640 1880 -620
rect 1900 -640 1920 -620
rect 1940 -640 1960 -620
rect 1980 -640 2000 -620
rect 2020 -640 2040 -620
rect 2060 -640 2080 -620
rect 2100 -640 2120 -620
rect 2140 -640 2160 -620
rect 2180 -640 2200 -620
rect 2220 -640 2240 -620
rect 2260 -640 2280 -620
rect 2300 -640 2320 -620
rect 2340 -640 2360 -620
rect 2380 -640 2400 -620
rect 2420 -640 2440 -620
rect 2460 -640 2480 -620
rect 2500 -640 2520 -620
rect 2540 -640 2560 -620
rect 2590 -640 2605 -620
rect 105 -655 2605 -640
rect 105 -715 2605 -700
rect 105 -735 120 -715
rect 140 -735 160 -715
rect 180 -735 200 -715
rect 220 -735 240 -715
rect 260 -735 280 -715
rect 300 -735 320 -715
rect 340 -735 360 -715
rect 380 -735 400 -715
rect 420 -735 440 -715
rect 460 -735 480 -715
rect 500 -735 520 -715
rect 540 -735 560 -715
rect 580 -735 600 -715
rect 620 -735 640 -715
rect 660 -735 680 -715
rect 700 -735 720 -715
rect 740 -735 760 -715
rect 780 -735 800 -715
rect 820 -735 840 -715
rect 860 -735 880 -715
rect 900 -735 920 -715
rect 940 -735 960 -715
rect 980 -735 1000 -715
rect 1020 -735 1040 -715
rect 1060 -735 1080 -715
rect 1100 -735 1120 -715
rect 1140 -735 1160 -715
rect 1180 -735 1200 -715
rect 1220 -735 1240 -715
rect 1260 -735 1280 -715
rect 1300 -735 1320 -715
rect 1340 -735 1360 -715
rect 1380 -735 1400 -715
rect 1420 -735 1440 -715
rect 1460 -735 1480 -715
rect 1500 -735 1520 -715
rect 1540 -735 1560 -715
rect 1580 -735 1600 -715
rect 1620 -735 1640 -715
rect 1660 -735 1680 -715
rect 1700 -735 1720 -715
rect 1740 -735 1760 -715
rect 1780 -735 1800 -715
rect 1820 -735 1840 -715
rect 1860 -735 1880 -715
rect 1900 -735 1920 -715
rect 1940 -735 1960 -715
rect 1980 -735 2000 -715
rect 2020 -735 2040 -715
rect 2060 -735 2080 -715
rect 2100 -735 2120 -715
rect 2140 -735 2160 -715
rect 2180 -735 2200 -715
rect 2220 -735 2240 -715
rect 2260 -735 2280 -715
rect 2300 -735 2320 -715
rect 2340 -735 2360 -715
rect 2380 -735 2400 -715
rect 2420 -735 2440 -715
rect 2460 -735 2480 -715
rect 2500 -735 2520 -715
rect 2540 -735 2560 -715
rect 2590 -735 2605 -715
rect 105 -750 2605 -735
rect 105 -810 2605 -795
rect 105 -830 120 -810
rect 140 -830 160 -810
rect 180 -830 200 -810
rect 220 -830 240 -810
rect 260 -830 280 -810
rect 300 -830 320 -810
rect 340 -830 360 -810
rect 380 -830 400 -810
rect 420 -830 440 -810
rect 460 -830 480 -810
rect 500 -830 520 -810
rect 540 -830 560 -810
rect 580 -830 600 -810
rect 620 -830 640 -810
rect 660 -830 680 -810
rect 700 -830 720 -810
rect 740 -830 760 -810
rect 780 -830 800 -810
rect 820 -830 840 -810
rect 860 -830 880 -810
rect 900 -830 920 -810
rect 940 -830 960 -810
rect 980 -830 1000 -810
rect 1020 -830 1040 -810
rect 1060 -830 1080 -810
rect 1100 -830 1120 -810
rect 1140 -830 1160 -810
rect 1180 -830 1200 -810
rect 1220 -830 1240 -810
rect 1260 -830 1280 -810
rect 1300 -830 1320 -810
rect 1340 -830 1360 -810
rect 1380 -830 1400 -810
rect 1420 -830 1440 -810
rect 1460 -830 1480 -810
rect 1500 -830 1520 -810
rect 1540 -830 1560 -810
rect 1580 -830 1600 -810
rect 1620 -830 1640 -810
rect 1660 -830 1680 -810
rect 1700 -830 1720 -810
rect 1740 -830 1760 -810
rect 1780 -830 1800 -810
rect 1820 -830 1840 -810
rect 1860 -830 1880 -810
rect 1900 -830 1920 -810
rect 1940 -830 1960 -810
rect 1980 -830 2000 -810
rect 2020 -830 2040 -810
rect 2060 -830 2080 -810
rect 2100 -830 2120 -810
rect 2140 -830 2160 -810
rect 2180 -830 2200 -810
rect 2220 -830 2240 -810
rect 2260 -830 2280 -810
rect 2300 -830 2320 -810
rect 2340 -830 2360 -810
rect 2380 -830 2400 -810
rect 2420 -830 2440 -810
rect 2460 -830 2480 -810
rect 2500 -830 2520 -810
rect 2540 -830 2560 -810
rect 2590 -830 2605 -810
rect 105 -845 2605 -830
rect 105 -905 2605 -890
rect 105 -925 120 -905
rect 140 -925 160 -905
rect 180 -925 200 -905
rect 220 -925 240 -905
rect 260 -925 280 -905
rect 300 -925 320 -905
rect 340 -925 360 -905
rect 380 -925 400 -905
rect 420 -925 440 -905
rect 460 -925 480 -905
rect 500 -925 520 -905
rect 540 -925 560 -905
rect 580 -925 600 -905
rect 620 -925 640 -905
rect 660 -925 680 -905
rect 700 -925 720 -905
rect 740 -925 760 -905
rect 780 -925 800 -905
rect 820 -925 840 -905
rect 860 -925 880 -905
rect 900 -925 920 -905
rect 940 -925 960 -905
rect 980 -925 1000 -905
rect 1020 -925 1040 -905
rect 1060 -925 1080 -905
rect 1100 -925 1120 -905
rect 1140 -925 1160 -905
rect 1180 -925 1200 -905
rect 1220 -925 1240 -905
rect 1260 -925 1280 -905
rect 1300 -925 1320 -905
rect 1340 -925 1360 -905
rect 1380 -925 1400 -905
rect 1420 -925 1440 -905
rect 1460 -925 1480 -905
rect 1500 -925 1520 -905
rect 1540 -925 1560 -905
rect 1580 -925 1600 -905
rect 1620 -925 1640 -905
rect 1660 -925 1680 -905
rect 1700 -925 1720 -905
rect 1740 -925 1760 -905
rect 1780 -925 1800 -905
rect 1820 -925 1840 -905
rect 1860 -925 1880 -905
rect 1900 -925 1920 -905
rect 1940 -925 1960 -905
rect 1980 -925 2000 -905
rect 2020 -925 2040 -905
rect 2060 -925 2080 -905
rect 2100 -925 2120 -905
rect 2140 -925 2160 -905
rect 2180 -925 2200 -905
rect 2220 -925 2240 -905
rect 2260 -925 2280 -905
rect 2300 -925 2320 -905
rect 2340 -925 2360 -905
rect 2380 -925 2400 -905
rect 2420 -925 2440 -905
rect 2460 -925 2480 -905
rect 2500 -925 2520 -905
rect 2540 -925 2560 -905
rect 2590 -925 2605 -905
rect 105 -940 2605 -925
rect 105 -1000 2605 -985
rect 105 -1020 120 -1000
rect 140 -1020 160 -1000
rect 180 -1020 200 -1000
rect 220 -1020 240 -1000
rect 260 -1020 280 -1000
rect 300 -1020 320 -1000
rect 340 -1020 360 -1000
rect 380 -1020 400 -1000
rect 420 -1020 440 -1000
rect 460 -1020 480 -1000
rect 500 -1020 520 -1000
rect 540 -1020 560 -1000
rect 580 -1020 600 -1000
rect 620 -1020 640 -1000
rect 660 -1020 680 -1000
rect 700 -1020 720 -1000
rect 740 -1020 760 -1000
rect 780 -1020 800 -1000
rect 820 -1020 840 -1000
rect 860 -1020 880 -1000
rect 900 -1020 920 -1000
rect 940 -1020 960 -1000
rect 980 -1020 1000 -1000
rect 1020 -1020 1040 -1000
rect 1060 -1020 1080 -1000
rect 1100 -1020 1120 -1000
rect 1140 -1020 1160 -1000
rect 1180 -1020 1200 -1000
rect 1220 -1020 1240 -1000
rect 1260 -1020 1280 -1000
rect 1300 -1020 1320 -1000
rect 1340 -1020 1360 -1000
rect 1380 -1020 1400 -1000
rect 1420 -1020 1440 -1000
rect 1460 -1020 1480 -1000
rect 1500 -1020 1520 -1000
rect 1540 -1020 1560 -1000
rect 1580 -1020 1600 -1000
rect 1620 -1020 1640 -1000
rect 1660 -1020 1680 -1000
rect 1700 -1020 1720 -1000
rect 1740 -1020 1760 -1000
rect 1780 -1020 1800 -1000
rect 1820 -1020 1840 -1000
rect 1860 -1020 1880 -1000
rect 1900 -1020 1920 -1000
rect 1940 -1020 1960 -1000
rect 1980 -1020 2000 -1000
rect 2020 -1020 2040 -1000
rect 2060 -1020 2080 -1000
rect 2100 -1020 2120 -1000
rect 2140 -1020 2160 -1000
rect 2180 -1020 2200 -1000
rect 2220 -1020 2240 -1000
rect 2260 -1020 2280 -1000
rect 2300 -1020 2320 -1000
rect 2340 -1020 2360 -1000
rect 2380 -1020 2400 -1000
rect 2420 -1020 2440 -1000
rect 2460 -1020 2480 -1000
rect 2500 -1020 2520 -1000
rect 2540 -1020 2560 -1000
rect 2590 -1020 2605 -1000
rect 105 -1035 2605 -1020
rect 105 -1095 2605 -1080
rect 105 -1115 120 -1095
rect 140 -1115 160 -1095
rect 180 -1115 200 -1095
rect 220 -1115 240 -1095
rect 260 -1115 280 -1095
rect 300 -1115 320 -1095
rect 340 -1115 360 -1095
rect 380 -1115 400 -1095
rect 420 -1115 440 -1095
rect 460 -1115 480 -1095
rect 500 -1115 520 -1095
rect 540 -1115 560 -1095
rect 580 -1115 600 -1095
rect 620 -1115 640 -1095
rect 660 -1115 680 -1095
rect 700 -1115 720 -1095
rect 740 -1115 760 -1095
rect 780 -1115 800 -1095
rect 820 -1115 840 -1095
rect 860 -1115 880 -1095
rect 900 -1115 920 -1095
rect 940 -1115 960 -1095
rect 980 -1115 1000 -1095
rect 1020 -1115 1040 -1095
rect 1060 -1115 1080 -1095
rect 1100 -1115 1120 -1095
rect 1140 -1115 1160 -1095
rect 1180 -1115 1200 -1095
rect 1220 -1115 1240 -1095
rect 1260 -1115 1280 -1095
rect 1300 -1115 1320 -1095
rect 1340 -1115 1360 -1095
rect 1380 -1115 1400 -1095
rect 1420 -1115 1440 -1095
rect 1460 -1115 1480 -1095
rect 1500 -1115 1520 -1095
rect 1540 -1115 1560 -1095
rect 1580 -1115 1600 -1095
rect 1620 -1115 1640 -1095
rect 1660 -1115 1680 -1095
rect 1700 -1115 1720 -1095
rect 1740 -1115 1760 -1095
rect 1780 -1115 1800 -1095
rect 1820 -1115 1840 -1095
rect 1860 -1115 1880 -1095
rect 1900 -1115 1920 -1095
rect 1940 -1115 1960 -1095
rect 1980 -1115 2000 -1095
rect 2020 -1115 2040 -1095
rect 2060 -1115 2080 -1095
rect 2100 -1115 2120 -1095
rect 2140 -1115 2160 -1095
rect 2180 -1115 2200 -1095
rect 2220 -1115 2240 -1095
rect 2260 -1115 2280 -1095
rect 2300 -1115 2320 -1095
rect 2340 -1115 2360 -1095
rect 2380 -1115 2400 -1095
rect 2420 -1115 2440 -1095
rect 2460 -1115 2480 -1095
rect 2500 -1115 2520 -1095
rect 2540 -1115 2560 -1095
rect 2590 -1115 2605 -1095
rect 105 -1130 2605 -1115
rect 105 -1190 2605 -1175
rect 105 -1210 120 -1190
rect 140 -1210 160 -1190
rect 180 -1210 200 -1190
rect 220 -1210 240 -1190
rect 260 -1210 280 -1190
rect 300 -1210 320 -1190
rect 340 -1210 360 -1190
rect 380 -1210 400 -1190
rect 420 -1210 440 -1190
rect 460 -1210 480 -1190
rect 500 -1210 520 -1190
rect 540 -1210 560 -1190
rect 580 -1210 600 -1190
rect 620 -1210 640 -1190
rect 660 -1210 680 -1190
rect 700 -1210 720 -1190
rect 740 -1210 760 -1190
rect 780 -1210 800 -1190
rect 820 -1210 840 -1190
rect 860 -1210 880 -1190
rect 900 -1210 920 -1190
rect 940 -1210 960 -1190
rect 980 -1210 1000 -1190
rect 1020 -1210 1040 -1190
rect 1060 -1210 1080 -1190
rect 1100 -1210 1120 -1190
rect 1140 -1210 1160 -1190
rect 1180 -1210 1200 -1190
rect 1220 -1210 1240 -1190
rect 1260 -1210 1280 -1190
rect 1300 -1210 1320 -1190
rect 1340 -1210 1360 -1190
rect 1380 -1210 1400 -1190
rect 1420 -1210 1440 -1190
rect 1460 -1210 1480 -1190
rect 1500 -1210 1520 -1190
rect 1540 -1210 1560 -1190
rect 1580 -1210 1600 -1190
rect 1620 -1210 1640 -1190
rect 1660 -1210 1680 -1190
rect 1700 -1210 1720 -1190
rect 1740 -1210 1760 -1190
rect 1780 -1210 1800 -1190
rect 1820 -1210 1840 -1190
rect 1860 -1210 1880 -1190
rect 1900 -1210 1920 -1190
rect 1940 -1210 1960 -1190
rect 1980 -1210 2000 -1190
rect 2020 -1210 2040 -1190
rect 2060 -1210 2080 -1190
rect 2100 -1210 2120 -1190
rect 2140 -1210 2160 -1190
rect 2180 -1210 2200 -1190
rect 2220 -1210 2240 -1190
rect 2260 -1210 2280 -1190
rect 2300 -1210 2320 -1190
rect 2340 -1210 2360 -1190
rect 2380 -1210 2400 -1190
rect 2420 -1210 2440 -1190
rect 2460 -1210 2480 -1190
rect 2500 -1210 2520 -1190
rect 2540 -1210 2560 -1190
rect 2590 -1210 2605 -1190
rect 105 -1225 2605 -1210
rect 105 -1285 2605 -1270
rect 105 -1305 120 -1285
rect 140 -1305 160 -1285
rect 180 -1305 200 -1285
rect 220 -1305 240 -1285
rect 260 -1305 280 -1285
rect 300 -1305 320 -1285
rect 340 -1305 360 -1285
rect 380 -1305 400 -1285
rect 420 -1305 440 -1285
rect 460 -1305 480 -1285
rect 500 -1305 520 -1285
rect 540 -1305 560 -1285
rect 580 -1305 600 -1285
rect 620 -1305 640 -1285
rect 660 -1305 680 -1285
rect 700 -1305 720 -1285
rect 740 -1305 760 -1285
rect 780 -1305 800 -1285
rect 820 -1305 840 -1285
rect 860 -1305 880 -1285
rect 900 -1305 920 -1285
rect 940 -1305 960 -1285
rect 980 -1305 1000 -1285
rect 1020 -1305 1040 -1285
rect 1060 -1305 1080 -1285
rect 1100 -1305 1120 -1285
rect 1140 -1305 1160 -1285
rect 1180 -1305 1200 -1285
rect 1220 -1305 1240 -1285
rect 1260 -1305 1280 -1285
rect 1300 -1305 1320 -1285
rect 1340 -1305 1360 -1285
rect 1380 -1305 1400 -1285
rect 1420 -1305 1440 -1285
rect 1460 -1305 1480 -1285
rect 1500 -1305 1520 -1285
rect 1540 -1305 1560 -1285
rect 1580 -1305 1600 -1285
rect 1620 -1305 1640 -1285
rect 1660 -1305 1680 -1285
rect 1700 -1305 1720 -1285
rect 1740 -1305 1760 -1285
rect 1780 -1305 1800 -1285
rect 1820 -1305 1840 -1285
rect 1860 -1305 1880 -1285
rect 1900 -1305 1920 -1285
rect 1940 -1305 1960 -1285
rect 1980 -1305 2000 -1285
rect 2020 -1305 2040 -1285
rect 2060 -1305 2080 -1285
rect 2100 -1305 2120 -1285
rect 2140 -1305 2160 -1285
rect 2180 -1305 2200 -1285
rect 2220 -1305 2240 -1285
rect 2260 -1305 2280 -1285
rect 2300 -1305 2320 -1285
rect 2340 -1305 2360 -1285
rect 2380 -1305 2400 -1285
rect 2420 -1305 2440 -1285
rect 2460 -1305 2480 -1285
rect 2500 -1305 2520 -1285
rect 2540 -1305 2560 -1285
rect 2590 -1305 2605 -1285
rect 105 -1320 2605 -1305
rect 105 -1380 2605 -1365
rect 105 -1400 120 -1380
rect 140 -1400 160 -1380
rect 180 -1400 200 -1380
rect 220 -1400 240 -1380
rect 260 -1400 280 -1380
rect 300 -1400 320 -1380
rect 340 -1400 360 -1380
rect 380 -1400 400 -1380
rect 420 -1400 440 -1380
rect 460 -1400 480 -1380
rect 500 -1400 520 -1380
rect 540 -1400 560 -1380
rect 580 -1400 600 -1380
rect 620 -1400 640 -1380
rect 660 -1400 680 -1380
rect 700 -1400 720 -1380
rect 740 -1400 760 -1380
rect 780 -1400 800 -1380
rect 820 -1400 840 -1380
rect 860 -1400 880 -1380
rect 900 -1400 920 -1380
rect 940 -1400 960 -1380
rect 980 -1400 1000 -1380
rect 1020 -1400 1040 -1380
rect 1060 -1400 1080 -1380
rect 1100 -1400 1120 -1380
rect 1140 -1400 1160 -1380
rect 1180 -1400 1200 -1380
rect 1220 -1400 1240 -1380
rect 1260 -1400 1280 -1380
rect 1300 -1400 1320 -1380
rect 1340 -1400 1360 -1380
rect 1380 -1400 1400 -1380
rect 1420 -1400 1440 -1380
rect 1460 -1400 1480 -1380
rect 1500 -1400 1520 -1380
rect 1540 -1400 1560 -1380
rect 1580 -1400 1600 -1380
rect 1620 -1400 1640 -1380
rect 1660 -1400 1680 -1380
rect 1700 -1400 1720 -1380
rect 1740 -1400 1760 -1380
rect 1780 -1400 1800 -1380
rect 1820 -1400 1840 -1380
rect 1860 -1400 1880 -1380
rect 1900 -1400 1920 -1380
rect 1940 -1400 1960 -1380
rect 1980 -1400 2000 -1380
rect 2020 -1400 2040 -1380
rect 2060 -1400 2080 -1380
rect 2100 -1400 2120 -1380
rect 2140 -1400 2160 -1380
rect 2180 -1400 2200 -1380
rect 2220 -1400 2240 -1380
rect 2260 -1400 2280 -1380
rect 2300 -1400 2320 -1380
rect 2340 -1400 2360 -1380
rect 2380 -1400 2400 -1380
rect 2420 -1400 2440 -1380
rect 2460 -1400 2480 -1380
rect 2500 -1400 2520 -1380
rect 2540 -1400 2560 -1380
rect 2590 -1400 2605 -1380
rect 105 -1415 2605 -1400
rect 105 -1475 2605 -1460
rect 105 -1495 120 -1475
rect 140 -1495 160 -1475
rect 180 -1495 200 -1475
rect 220 -1495 240 -1475
rect 260 -1495 280 -1475
rect 300 -1495 320 -1475
rect 340 -1495 360 -1475
rect 380 -1495 400 -1475
rect 420 -1495 440 -1475
rect 460 -1495 480 -1475
rect 500 -1495 520 -1475
rect 540 -1495 560 -1475
rect 580 -1495 600 -1475
rect 620 -1495 640 -1475
rect 660 -1495 680 -1475
rect 700 -1495 720 -1475
rect 740 -1495 760 -1475
rect 780 -1495 800 -1475
rect 820 -1495 840 -1475
rect 860 -1495 880 -1475
rect 900 -1495 920 -1475
rect 940 -1495 960 -1475
rect 980 -1495 1000 -1475
rect 1020 -1495 1040 -1475
rect 1060 -1495 1080 -1475
rect 1100 -1495 1120 -1475
rect 1140 -1495 1160 -1475
rect 1180 -1495 1200 -1475
rect 1220 -1495 1240 -1475
rect 1260 -1495 1280 -1475
rect 1300 -1495 1320 -1475
rect 1340 -1495 1360 -1475
rect 1380 -1495 1400 -1475
rect 1420 -1495 1440 -1475
rect 1460 -1495 1480 -1475
rect 1500 -1495 1520 -1475
rect 1540 -1495 1560 -1475
rect 1580 -1495 1600 -1475
rect 1620 -1495 1640 -1475
rect 1660 -1495 1680 -1475
rect 1700 -1495 1720 -1475
rect 1740 -1495 1760 -1475
rect 1780 -1495 1800 -1475
rect 1820 -1495 1840 -1475
rect 1860 -1495 1880 -1475
rect 1900 -1495 1920 -1475
rect 1940 -1495 1960 -1475
rect 1980 -1495 2000 -1475
rect 2020 -1495 2040 -1475
rect 2060 -1495 2080 -1475
rect 2100 -1495 2120 -1475
rect 2140 -1495 2160 -1475
rect 2180 -1495 2200 -1475
rect 2220 -1495 2240 -1475
rect 2260 -1495 2280 -1475
rect 2300 -1495 2320 -1475
rect 2340 -1495 2360 -1475
rect 2380 -1495 2400 -1475
rect 2420 -1495 2440 -1475
rect 2460 -1495 2480 -1475
rect 2500 -1495 2520 -1475
rect 2540 -1495 2560 -1475
rect 2590 -1495 2605 -1475
rect 105 -1510 2605 -1495
rect 105 -1570 2605 -1555
rect 105 -1590 120 -1570
rect 140 -1590 160 -1570
rect 180 -1590 200 -1570
rect 220 -1590 240 -1570
rect 260 -1590 280 -1570
rect 300 -1590 320 -1570
rect 340 -1590 360 -1570
rect 380 -1590 400 -1570
rect 420 -1590 440 -1570
rect 460 -1590 480 -1570
rect 500 -1590 520 -1570
rect 540 -1590 560 -1570
rect 580 -1590 600 -1570
rect 620 -1590 640 -1570
rect 660 -1590 680 -1570
rect 700 -1590 720 -1570
rect 740 -1590 760 -1570
rect 780 -1590 800 -1570
rect 820 -1590 840 -1570
rect 860 -1590 880 -1570
rect 900 -1590 920 -1570
rect 940 -1590 960 -1570
rect 980 -1590 1000 -1570
rect 1020 -1590 1040 -1570
rect 1060 -1590 1080 -1570
rect 1100 -1590 1120 -1570
rect 1140 -1590 1160 -1570
rect 1180 -1590 1200 -1570
rect 1220 -1590 1240 -1570
rect 1260 -1590 1280 -1570
rect 1300 -1590 1320 -1570
rect 1340 -1590 1360 -1570
rect 1380 -1590 1400 -1570
rect 1420 -1590 1440 -1570
rect 1460 -1590 1480 -1570
rect 1500 -1590 1520 -1570
rect 1540 -1590 1560 -1570
rect 1580 -1590 1600 -1570
rect 1620 -1590 1640 -1570
rect 1660 -1590 1680 -1570
rect 1700 -1590 1720 -1570
rect 1740 -1590 1760 -1570
rect 1780 -1590 1800 -1570
rect 1820 -1590 1840 -1570
rect 1860 -1590 1880 -1570
rect 1900 -1590 1920 -1570
rect 1940 -1590 1960 -1570
rect 1980 -1590 2000 -1570
rect 2020 -1590 2040 -1570
rect 2060 -1590 2080 -1570
rect 2100 -1590 2120 -1570
rect 2140 -1590 2160 -1570
rect 2180 -1590 2200 -1570
rect 2220 -1590 2240 -1570
rect 2260 -1590 2280 -1570
rect 2300 -1590 2320 -1570
rect 2340 -1590 2360 -1570
rect 2380 -1590 2400 -1570
rect 2420 -1590 2440 -1570
rect 2460 -1590 2480 -1570
rect 2500 -1590 2520 -1570
rect 2540 -1590 2560 -1570
rect 2590 -1590 2605 -1570
rect 105 -1605 2605 -1590
rect 105 -1665 2605 -1650
rect 105 -1685 120 -1665
rect 140 -1685 160 -1665
rect 180 -1685 200 -1665
rect 220 -1685 240 -1665
rect 260 -1685 280 -1665
rect 300 -1685 320 -1665
rect 340 -1685 360 -1665
rect 380 -1685 400 -1665
rect 420 -1685 440 -1665
rect 460 -1685 480 -1665
rect 500 -1685 520 -1665
rect 540 -1685 560 -1665
rect 580 -1685 600 -1665
rect 620 -1685 640 -1665
rect 660 -1685 680 -1665
rect 700 -1685 720 -1665
rect 740 -1685 760 -1665
rect 780 -1685 800 -1665
rect 820 -1685 840 -1665
rect 860 -1685 880 -1665
rect 900 -1685 920 -1665
rect 940 -1685 960 -1665
rect 980 -1685 1000 -1665
rect 1020 -1685 1040 -1665
rect 1060 -1685 1080 -1665
rect 1100 -1685 1120 -1665
rect 1140 -1685 1160 -1665
rect 1180 -1685 1200 -1665
rect 1220 -1685 1240 -1665
rect 1260 -1685 1280 -1665
rect 1300 -1685 1320 -1665
rect 1340 -1685 1360 -1665
rect 1380 -1685 1400 -1665
rect 1420 -1685 1440 -1665
rect 1460 -1685 1480 -1665
rect 1500 -1685 1520 -1665
rect 1540 -1685 1560 -1665
rect 1580 -1685 1600 -1665
rect 1620 -1685 1640 -1665
rect 1660 -1685 1680 -1665
rect 1700 -1685 1720 -1665
rect 1740 -1685 1760 -1665
rect 1780 -1685 1800 -1665
rect 1820 -1685 1840 -1665
rect 1860 -1685 1880 -1665
rect 1900 -1685 1920 -1665
rect 1940 -1685 1960 -1665
rect 1980 -1685 2000 -1665
rect 2020 -1685 2040 -1665
rect 2060 -1685 2080 -1665
rect 2100 -1685 2120 -1665
rect 2140 -1685 2160 -1665
rect 2180 -1685 2200 -1665
rect 2220 -1685 2240 -1665
rect 2260 -1685 2280 -1665
rect 2300 -1685 2320 -1665
rect 2340 -1685 2360 -1665
rect 2380 -1685 2400 -1665
rect 2420 -1685 2440 -1665
rect 2460 -1685 2480 -1665
rect 2500 -1685 2520 -1665
rect 2540 -1685 2560 -1665
rect 2590 -1685 2605 -1665
rect 105 -1700 2605 -1685
rect 105 -1760 2605 -1745
rect 105 -1780 120 -1760
rect 140 -1780 160 -1760
rect 180 -1780 200 -1760
rect 220 -1780 240 -1760
rect 260 -1780 280 -1760
rect 300 -1780 320 -1760
rect 340 -1780 360 -1760
rect 380 -1780 400 -1760
rect 420 -1780 440 -1760
rect 460 -1780 480 -1760
rect 500 -1780 520 -1760
rect 540 -1780 560 -1760
rect 580 -1780 600 -1760
rect 620 -1780 640 -1760
rect 660 -1780 680 -1760
rect 700 -1780 720 -1760
rect 740 -1780 760 -1760
rect 780 -1780 800 -1760
rect 820 -1780 840 -1760
rect 860 -1780 880 -1760
rect 900 -1780 920 -1760
rect 940 -1780 960 -1760
rect 980 -1780 1000 -1760
rect 1020 -1780 1040 -1760
rect 1060 -1780 1080 -1760
rect 1100 -1780 1120 -1760
rect 1140 -1780 1160 -1760
rect 1180 -1780 1200 -1760
rect 1220 -1780 1240 -1760
rect 1260 -1780 1280 -1760
rect 1300 -1780 1320 -1760
rect 1340 -1780 1360 -1760
rect 1380 -1780 1400 -1760
rect 1420 -1780 1440 -1760
rect 1460 -1780 1480 -1760
rect 1500 -1780 1520 -1760
rect 1540 -1780 1560 -1760
rect 1580 -1780 1600 -1760
rect 1620 -1780 1640 -1760
rect 1660 -1780 1680 -1760
rect 1700 -1780 1720 -1760
rect 1740 -1780 1760 -1760
rect 1780 -1780 1800 -1760
rect 1820 -1780 1840 -1760
rect 1860 -1780 1880 -1760
rect 1900 -1780 1920 -1760
rect 1940 -1780 1960 -1760
rect 1980 -1780 2000 -1760
rect 2020 -1780 2040 -1760
rect 2060 -1780 2080 -1760
rect 2100 -1780 2120 -1760
rect 2140 -1780 2160 -1760
rect 2180 -1780 2200 -1760
rect 2220 -1780 2240 -1760
rect 2260 -1780 2280 -1760
rect 2300 -1780 2320 -1760
rect 2340 -1780 2360 -1760
rect 2380 -1780 2400 -1760
rect 2420 -1780 2440 -1760
rect 2460 -1780 2480 -1760
rect 2500 -1780 2520 -1760
rect 2540 -1780 2560 -1760
rect 2590 -1780 2605 -1760
rect 105 -1795 2605 -1780
rect 105 -1855 2605 -1840
rect 105 -1875 120 -1855
rect 140 -1875 160 -1855
rect 180 -1875 200 -1855
rect 220 -1875 240 -1855
rect 260 -1875 280 -1855
rect 300 -1875 320 -1855
rect 340 -1875 360 -1855
rect 380 -1875 400 -1855
rect 420 -1875 440 -1855
rect 460 -1875 480 -1855
rect 500 -1875 520 -1855
rect 540 -1875 560 -1855
rect 580 -1875 600 -1855
rect 620 -1875 640 -1855
rect 660 -1875 680 -1855
rect 700 -1875 720 -1855
rect 740 -1875 760 -1855
rect 780 -1875 800 -1855
rect 820 -1875 840 -1855
rect 860 -1875 880 -1855
rect 900 -1875 920 -1855
rect 940 -1875 960 -1855
rect 980 -1875 1000 -1855
rect 1020 -1875 1040 -1855
rect 1060 -1875 1080 -1855
rect 1100 -1875 1120 -1855
rect 1140 -1875 1160 -1855
rect 1180 -1875 1200 -1855
rect 1220 -1875 1240 -1855
rect 1260 -1875 1280 -1855
rect 1300 -1875 1320 -1855
rect 1340 -1875 1360 -1855
rect 1380 -1875 1400 -1855
rect 1420 -1875 1440 -1855
rect 1460 -1875 1480 -1855
rect 1500 -1875 1520 -1855
rect 1540 -1875 1560 -1855
rect 1580 -1875 1600 -1855
rect 1620 -1875 1640 -1855
rect 1660 -1875 1680 -1855
rect 1700 -1875 1720 -1855
rect 1740 -1875 1760 -1855
rect 1780 -1875 1800 -1855
rect 1820 -1875 1840 -1855
rect 1860 -1875 1880 -1855
rect 1900 -1875 1920 -1855
rect 1940 -1875 1960 -1855
rect 1980 -1875 2000 -1855
rect 2020 -1875 2040 -1855
rect 2060 -1875 2080 -1855
rect 2100 -1875 2120 -1855
rect 2140 -1875 2160 -1855
rect 2180 -1875 2200 -1855
rect 2220 -1875 2240 -1855
rect 2260 -1875 2280 -1855
rect 2300 -1875 2320 -1855
rect 2340 -1875 2360 -1855
rect 2380 -1875 2400 -1855
rect 2420 -1875 2440 -1855
rect 2460 -1875 2480 -1855
rect 2500 -1875 2520 -1855
rect 2540 -1875 2560 -1855
rect 2590 -1875 2605 -1855
rect 105 -1890 2605 -1875
rect 105 -1950 2605 -1935
rect 105 -1970 120 -1950
rect 140 -1970 160 -1950
rect 180 -1970 200 -1950
rect 220 -1970 240 -1950
rect 260 -1970 280 -1950
rect 300 -1970 320 -1950
rect 340 -1970 360 -1950
rect 380 -1970 400 -1950
rect 420 -1970 440 -1950
rect 460 -1970 480 -1950
rect 500 -1970 520 -1950
rect 540 -1970 560 -1950
rect 580 -1970 600 -1950
rect 620 -1970 640 -1950
rect 660 -1970 680 -1950
rect 700 -1970 720 -1950
rect 740 -1970 760 -1950
rect 780 -1970 800 -1950
rect 820 -1970 840 -1950
rect 860 -1970 880 -1950
rect 900 -1970 920 -1950
rect 940 -1970 960 -1950
rect 980 -1970 1000 -1950
rect 1020 -1970 1040 -1950
rect 1060 -1970 1080 -1950
rect 1100 -1970 1120 -1950
rect 1140 -1970 1160 -1950
rect 1180 -1970 1200 -1950
rect 1220 -1970 1240 -1950
rect 1260 -1970 1280 -1950
rect 1300 -1970 1320 -1950
rect 1340 -1970 1360 -1950
rect 1380 -1970 1400 -1950
rect 1420 -1970 1440 -1950
rect 1460 -1970 1480 -1950
rect 1500 -1970 1520 -1950
rect 1540 -1970 1560 -1950
rect 1580 -1970 1600 -1950
rect 1620 -1970 1640 -1950
rect 1660 -1970 1680 -1950
rect 1700 -1970 1720 -1950
rect 1740 -1970 1760 -1950
rect 1780 -1970 1800 -1950
rect 1820 -1970 1840 -1950
rect 1860 -1970 1880 -1950
rect 1900 -1970 1920 -1950
rect 1940 -1970 1960 -1950
rect 1980 -1970 2000 -1950
rect 2020 -1970 2040 -1950
rect 2060 -1970 2080 -1950
rect 2100 -1970 2120 -1950
rect 2140 -1970 2160 -1950
rect 2180 -1970 2200 -1950
rect 2220 -1970 2240 -1950
rect 2260 -1970 2280 -1950
rect 2300 -1970 2320 -1950
rect 2340 -1970 2360 -1950
rect 2380 -1970 2400 -1950
rect 2420 -1970 2440 -1950
rect 2460 -1970 2480 -1950
rect 2500 -1970 2520 -1950
rect 2540 -1970 2560 -1950
rect 2590 -1970 2605 -1950
rect 105 -1985 2605 -1970
rect 105 -2045 2605 -2030
rect 105 -2065 120 -2045
rect 140 -2065 160 -2045
rect 180 -2065 200 -2045
rect 220 -2065 240 -2045
rect 260 -2065 280 -2045
rect 300 -2065 320 -2045
rect 340 -2065 360 -2045
rect 380 -2065 400 -2045
rect 420 -2065 440 -2045
rect 460 -2065 480 -2045
rect 500 -2065 520 -2045
rect 540 -2065 560 -2045
rect 580 -2065 600 -2045
rect 620 -2065 640 -2045
rect 660 -2065 680 -2045
rect 700 -2065 720 -2045
rect 740 -2065 760 -2045
rect 780 -2065 800 -2045
rect 820 -2065 840 -2045
rect 860 -2065 880 -2045
rect 900 -2065 920 -2045
rect 940 -2065 960 -2045
rect 980 -2065 1000 -2045
rect 1020 -2065 1040 -2045
rect 1060 -2065 1080 -2045
rect 1100 -2065 1120 -2045
rect 1140 -2065 1160 -2045
rect 1180 -2065 1200 -2045
rect 1220 -2065 1240 -2045
rect 1260 -2065 1280 -2045
rect 1300 -2065 1320 -2045
rect 1340 -2065 1360 -2045
rect 1380 -2065 1400 -2045
rect 1420 -2065 1440 -2045
rect 1460 -2065 1480 -2045
rect 1500 -2065 1520 -2045
rect 1540 -2065 1560 -2045
rect 1580 -2065 1600 -2045
rect 1620 -2065 1640 -2045
rect 1660 -2065 1680 -2045
rect 1700 -2065 1720 -2045
rect 1740 -2065 1760 -2045
rect 1780 -2065 1800 -2045
rect 1820 -2065 1840 -2045
rect 1860 -2065 1880 -2045
rect 1900 -2065 1920 -2045
rect 1940 -2065 1960 -2045
rect 1980 -2065 2000 -2045
rect 2020 -2065 2040 -2045
rect 2060 -2065 2080 -2045
rect 2100 -2065 2120 -2045
rect 2140 -2065 2160 -2045
rect 2180 -2065 2200 -2045
rect 2220 -2065 2240 -2045
rect 2260 -2065 2280 -2045
rect 2300 -2065 2320 -2045
rect 2340 -2065 2360 -2045
rect 2380 -2065 2400 -2045
rect 2420 -2065 2440 -2045
rect 2460 -2065 2480 -2045
rect 2500 -2065 2520 -2045
rect 2540 -2065 2560 -2045
rect 2590 -2065 2605 -2045
rect 105 -2080 2605 -2065
rect 105 -2140 2605 -2125
rect 105 -2160 120 -2140
rect 140 -2160 160 -2140
rect 180 -2160 200 -2140
rect 220 -2160 240 -2140
rect 260 -2160 280 -2140
rect 300 -2160 320 -2140
rect 340 -2160 360 -2140
rect 380 -2160 400 -2140
rect 420 -2160 440 -2140
rect 460 -2160 480 -2140
rect 500 -2160 520 -2140
rect 540 -2160 560 -2140
rect 580 -2160 600 -2140
rect 620 -2160 640 -2140
rect 660 -2160 680 -2140
rect 700 -2160 720 -2140
rect 740 -2160 760 -2140
rect 780 -2160 800 -2140
rect 820 -2160 840 -2140
rect 860 -2160 880 -2140
rect 900 -2160 920 -2140
rect 940 -2160 960 -2140
rect 980 -2160 1000 -2140
rect 1020 -2160 1040 -2140
rect 1060 -2160 1080 -2140
rect 1100 -2160 1120 -2140
rect 1140 -2160 1160 -2140
rect 1180 -2160 1200 -2140
rect 1220 -2160 1240 -2140
rect 1260 -2160 1280 -2140
rect 1300 -2160 1320 -2140
rect 1340 -2160 1360 -2140
rect 1380 -2160 1400 -2140
rect 1420 -2160 1440 -2140
rect 1460 -2160 1480 -2140
rect 1500 -2160 1520 -2140
rect 1540 -2160 1560 -2140
rect 1580 -2160 1600 -2140
rect 1620 -2160 1640 -2140
rect 1660 -2160 1680 -2140
rect 1700 -2160 1720 -2140
rect 1740 -2160 1760 -2140
rect 1780 -2160 1800 -2140
rect 1820 -2160 1840 -2140
rect 1860 -2160 1880 -2140
rect 1900 -2160 1920 -2140
rect 1940 -2160 1960 -2140
rect 1980 -2160 2000 -2140
rect 2020 -2160 2040 -2140
rect 2060 -2160 2080 -2140
rect 2100 -2160 2120 -2140
rect 2140 -2160 2160 -2140
rect 2180 -2160 2200 -2140
rect 2220 -2160 2240 -2140
rect 2260 -2160 2280 -2140
rect 2300 -2160 2320 -2140
rect 2340 -2160 2360 -2140
rect 2380 -2160 2400 -2140
rect 2420 -2160 2440 -2140
rect 2460 -2160 2480 -2140
rect 2500 -2160 2520 -2140
rect 2540 -2160 2560 -2140
rect 2590 -2160 2605 -2140
rect 105 -2175 2605 -2160
rect 105 -2235 2605 -2220
rect 105 -2255 120 -2235
rect 140 -2255 160 -2235
rect 180 -2255 200 -2235
rect 220 -2255 240 -2235
rect 260 -2255 280 -2235
rect 300 -2255 320 -2235
rect 340 -2255 360 -2235
rect 380 -2255 400 -2235
rect 420 -2255 440 -2235
rect 460 -2255 480 -2235
rect 500 -2255 520 -2235
rect 540 -2255 560 -2235
rect 580 -2255 600 -2235
rect 620 -2255 640 -2235
rect 660 -2255 680 -2235
rect 700 -2255 720 -2235
rect 740 -2255 760 -2235
rect 780 -2255 800 -2235
rect 820 -2255 840 -2235
rect 860 -2255 880 -2235
rect 900 -2255 920 -2235
rect 940 -2255 960 -2235
rect 980 -2255 1000 -2235
rect 1020 -2255 1040 -2235
rect 1060 -2255 1080 -2235
rect 1100 -2255 1120 -2235
rect 1140 -2255 1160 -2235
rect 1180 -2255 1200 -2235
rect 1220 -2255 1240 -2235
rect 1260 -2255 1280 -2235
rect 1300 -2255 1320 -2235
rect 1340 -2255 1360 -2235
rect 1380 -2255 1400 -2235
rect 1420 -2255 1440 -2235
rect 1460 -2255 1480 -2235
rect 1500 -2255 1520 -2235
rect 1540 -2255 1560 -2235
rect 1580 -2255 1600 -2235
rect 1620 -2255 1640 -2235
rect 1660 -2255 1680 -2235
rect 1700 -2255 1720 -2235
rect 1740 -2255 1760 -2235
rect 1780 -2255 1800 -2235
rect 1820 -2255 1840 -2235
rect 1860 -2255 1880 -2235
rect 1900 -2255 1920 -2235
rect 1940 -2255 1960 -2235
rect 1980 -2255 2000 -2235
rect 2020 -2255 2040 -2235
rect 2060 -2255 2080 -2235
rect 2100 -2255 2120 -2235
rect 2140 -2255 2160 -2235
rect 2180 -2255 2200 -2235
rect 2220 -2255 2240 -2235
rect 2260 -2255 2280 -2235
rect 2300 -2255 2320 -2235
rect 2340 -2255 2360 -2235
rect 2380 -2255 2400 -2235
rect 2420 -2255 2440 -2235
rect 2460 -2255 2480 -2235
rect 2500 -2255 2520 -2235
rect 2540 -2255 2560 -2235
rect 2590 -2255 2605 -2235
rect 105 -2270 2605 -2255
rect 105 -2330 2605 -2315
rect 105 -2350 120 -2330
rect 140 -2350 160 -2330
rect 180 -2350 200 -2330
rect 220 -2350 240 -2330
rect 260 -2350 280 -2330
rect 300 -2350 320 -2330
rect 340 -2350 360 -2330
rect 380 -2350 400 -2330
rect 420 -2350 440 -2330
rect 460 -2350 480 -2330
rect 500 -2350 520 -2330
rect 540 -2350 560 -2330
rect 580 -2350 600 -2330
rect 620 -2350 640 -2330
rect 660 -2350 680 -2330
rect 700 -2350 720 -2330
rect 740 -2350 760 -2330
rect 780 -2350 800 -2330
rect 820 -2350 840 -2330
rect 860 -2350 880 -2330
rect 900 -2350 920 -2330
rect 940 -2350 960 -2330
rect 980 -2350 1000 -2330
rect 1020 -2350 1040 -2330
rect 1060 -2350 1080 -2330
rect 1100 -2350 1120 -2330
rect 1140 -2350 1160 -2330
rect 1180 -2350 1200 -2330
rect 1220 -2350 1240 -2330
rect 1260 -2350 1280 -2330
rect 1300 -2350 1320 -2330
rect 1340 -2350 1360 -2330
rect 1380 -2350 1400 -2330
rect 1420 -2350 1440 -2330
rect 1460 -2350 1480 -2330
rect 1500 -2350 1520 -2330
rect 1540 -2350 1560 -2330
rect 1580 -2350 1600 -2330
rect 1620 -2350 1640 -2330
rect 1660 -2350 1680 -2330
rect 1700 -2350 1720 -2330
rect 1740 -2350 1760 -2330
rect 1780 -2350 1800 -2330
rect 1820 -2350 1840 -2330
rect 1860 -2350 1880 -2330
rect 1900 -2350 1920 -2330
rect 1940 -2350 1960 -2330
rect 1980 -2350 2000 -2330
rect 2020 -2350 2040 -2330
rect 2060 -2350 2080 -2330
rect 2100 -2350 2120 -2330
rect 2140 -2350 2160 -2330
rect 2180 -2350 2200 -2330
rect 2220 -2350 2240 -2330
rect 2260 -2350 2280 -2330
rect 2300 -2350 2320 -2330
rect 2340 -2350 2360 -2330
rect 2380 -2350 2400 -2330
rect 2420 -2350 2440 -2330
rect 2460 -2350 2480 -2330
rect 2500 -2350 2520 -2330
rect 2540 -2350 2560 -2330
rect 2590 -2350 2605 -2330
rect 105 -2365 2605 -2350
rect 105 -2425 2605 -2410
rect 105 -2445 120 -2425
rect 140 -2445 160 -2425
rect 180 -2445 200 -2425
rect 220 -2445 240 -2425
rect 260 -2445 280 -2425
rect 300 -2445 320 -2425
rect 340 -2445 360 -2425
rect 380 -2445 400 -2425
rect 420 -2445 440 -2425
rect 460 -2445 480 -2425
rect 500 -2445 520 -2425
rect 540 -2445 560 -2425
rect 580 -2445 600 -2425
rect 620 -2445 640 -2425
rect 660 -2445 680 -2425
rect 700 -2445 720 -2425
rect 740 -2445 760 -2425
rect 780 -2445 800 -2425
rect 820 -2445 840 -2425
rect 860 -2445 880 -2425
rect 900 -2445 920 -2425
rect 940 -2445 960 -2425
rect 980 -2445 1000 -2425
rect 1020 -2445 1040 -2425
rect 1060 -2445 1080 -2425
rect 1100 -2445 1120 -2425
rect 1140 -2445 1160 -2425
rect 1180 -2445 1200 -2425
rect 1220 -2445 1240 -2425
rect 1260 -2445 1280 -2425
rect 1300 -2445 1320 -2425
rect 1340 -2445 1360 -2425
rect 1380 -2445 1400 -2425
rect 1420 -2445 1440 -2425
rect 1460 -2445 1480 -2425
rect 1500 -2445 1520 -2425
rect 1540 -2445 1560 -2425
rect 1580 -2445 1600 -2425
rect 1620 -2445 1640 -2425
rect 1660 -2445 1680 -2425
rect 1700 -2445 1720 -2425
rect 1740 -2445 1760 -2425
rect 1780 -2445 1800 -2425
rect 1820 -2445 1840 -2425
rect 1860 -2445 1880 -2425
rect 1900 -2445 1920 -2425
rect 1940 -2445 1960 -2425
rect 1980 -2445 2000 -2425
rect 2020 -2445 2040 -2425
rect 2060 -2445 2080 -2425
rect 2100 -2445 2120 -2425
rect 2140 -2445 2160 -2425
rect 2180 -2445 2200 -2425
rect 2220 -2445 2240 -2425
rect 2260 -2445 2280 -2425
rect 2300 -2445 2320 -2425
rect 2340 -2445 2360 -2425
rect 2380 -2445 2400 -2425
rect 2420 -2445 2440 -2425
rect 2460 -2445 2480 -2425
rect 2500 -2445 2520 -2425
rect 2540 -2445 2560 -2425
rect 2590 -2445 2605 -2425
rect 105 -2460 2605 -2445
rect 105 -2520 2605 -2505
rect 105 -2540 120 -2520
rect 140 -2540 160 -2520
rect 180 -2540 200 -2520
rect 220 -2540 240 -2520
rect 260 -2540 280 -2520
rect 300 -2540 320 -2520
rect 340 -2540 360 -2520
rect 380 -2540 400 -2520
rect 420 -2540 440 -2520
rect 460 -2540 480 -2520
rect 500 -2540 520 -2520
rect 540 -2540 560 -2520
rect 580 -2540 600 -2520
rect 620 -2540 640 -2520
rect 660 -2540 680 -2520
rect 700 -2540 720 -2520
rect 740 -2540 760 -2520
rect 780 -2540 800 -2520
rect 820 -2540 840 -2520
rect 860 -2540 880 -2520
rect 900 -2540 920 -2520
rect 940 -2540 960 -2520
rect 980 -2540 1000 -2520
rect 1020 -2540 1040 -2520
rect 1060 -2540 1080 -2520
rect 1100 -2540 1120 -2520
rect 1140 -2540 1160 -2520
rect 1180 -2540 1200 -2520
rect 1220 -2540 1240 -2520
rect 1260 -2540 1280 -2520
rect 1300 -2540 1320 -2520
rect 1340 -2540 1360 -2520
rect 1380 -2540 1400 -2520
rect 1420 -2540 1440 -2520
rect 1460 -2540 1480 -2520
rect 1500 -2540 1520 -2520
rect 1540 -2540 1560 -2520
rect 1580 -2540 1600 -2520
rect 1620 -2540 1640 -2520
rect 1660 -2540 1680 -2520
rect 1700 -2540 1720 -2520
rect 1740 -2540 1760 -2520
rect 1780 -2540 1800 -2520
rect 1820 -2540 1840 -2520
rect 1860 -2540 1880 -2520
rect 1900 -2540 1920 -2520
rect 1940 -2540 1960 -2520
rect 1980 -2540 2000 -2520
rect 2020 -2540 2040 -2520
rect 2060 -2540 2080 -2520
rect 2100 -2540 2120 -2520
rect 2140 -2540 2160 -2520
rect 2180 -2540 2200 -2520
rect 2220 -2540 2240 -2520
rect 2260 -2540 2280 -2520
rect 2300 -2540 2320 -2520
rect 2340 -2540 2360 -2520
rect 2380 -2540 2400 -2520
rect 2420 -2540 2440 -2520
rect 2460 -2540 2480 -2520
rect 2500 -2540 2520 -2520
rect 2540 -2540 2560 -2520
rect 2590 -2540 2605 -2520
rect 105 -2550 2605 -2540
<< ndiffc >>
rect 200 2277 220 2297
rect 240 2277 260 2297
rect 280 2277 300 2297
rect 320 2277 340 2297
rect 360 2277 380 2297
rect 400 2277 420 2297
rect 440 2277 460 2297
rect 480 2277 500 2297
rect 520 2277 540 2297
rect 560 2277 580 2297
rect 600 2277 620 2297
rect 640 2277 660 2297
rect 680 2277 700 2297
rect 720 2277 740 2297
rect 760 2277 780 2297
rect 800 2277 820 2297
rect 840 2277 860 2297
rect 880 2277 900 2297
rect 920 2277 940 2297
rect 960 2277 980 2297
rect 1000 2277 1020 2297
rect 1040 2277 1060 2297
rect 1080 2277 1100 2297
rect 1120 2277 1140 2297
rect 1160 2277 1180 2297
rect 1200 2277 1220 2297
rect 1240 2277 1260 2297
rect 1280 2277 1300 2297
rect 1320 2277 1340 2297
rect 1360 2277 1380 2297
rect 1400 2277 1420 2297
rect 1440 2277 1460 2297
rect 1480 2277 1500 2297
rect 1520 2277 1540 2297
rect 1560 2277 1580 2297
rect 1600 2277 1620 2297
rect 1640 2277 1660 2297
rect 1680 2277 1700 2297
rect 1720 2277 1740 2297
rect 1760 2277 1780 2297
rect 1800 2277 1820 2297
rect 1840 2277 1860 2297
rect 1880 2277 1900 2297
rect 1920 2277 1940 2297
rect 1960 2277 1980 2297
rect 2000 2277 2020 2297
rect 2040 2277 2060 2297
rect 2080 2277 2100 2297
rect 2120 2277 2140 2297
rect 2160 2277 2180 2297
rect 2200 2277 2220 2297
rect 2240 2277 2260 2297
rect 2280 2277 2300 2297
rect 2320 2277 2340 2297
rect 2360 2277 2380 2297
rect 2400 2277 2420 2297
rect 2440 2277 2460 2297
rect 2480 2277 2500 2297
rect 2520 2277 2540 2297
rect 2560 2277 2580 2297
rect 2600 2277 2620 2297
rect 2640 2277 2660 2297
rect 200 2195 220 2215
rect 240 2195 260 2215
rect 280 2195 300 2215
rect 320 2195 340 2215
rect 360 2195 380 2215
rect 400 2195 420 2215
rect 440 2195 460 2215
rect 480 2195 500 2215
rect 520 2195 540 2215
rect 560 2195 580 2215
rect 600 2195 620 2215
rect 640 2195 660 2215
rect 680 2195 700 2215
rect 720 2195 740 2215
rect 760 2195 780 2215
rect 800 2195 820 2215
rect 840 2195 860 2215
rect 880 2195 900 2215
rect 920 2195 940 2215
rect 960 2195 980 2215
rect 1000 2195 1020 2215
rect 1040 2195 1060 2215
rect 1080 2195 1100 2215
rect 1120 2195 1140 2215
rect 1160 2195 1180 2215
rect 1200 2195 1220 2215
rect 1240 2195 1260 2215
rect 1280 2195 1300 2215
rect 1320 2195 1340 2215
rect 1360 2195 1380 2215
rect 1400 2195 1420 2215
rect 1440 2195 1460 2215
rect 1480 2195 1500 2215
rect 1520 2195 1540 2215
rect 1560 2195 1580 2215
rect 1600 2195 1620 2215
rect 1640 2195 1660 2215
rect 1680 2195 1700 2215
rect 1720 2195 1740 2215
rect 1760 2195 1780 2215
rect 1800 2195 1820 2215
rect 1840 2195 1860 2215
rect 1880 2195 1900 2215
rect 1920 2195 1940 2215
rect 1960 2195 1980 2215
rect 2000 2195 2020 2215
rect 2040 2195 2060 2215
rect 2080 2195 2100 2215
rect 2120 2195 2140 2215
rect 2160 2195 2180 2215
rect 2200 2195 2220 2215
rect 2240 2195 2260 2215
rect 2280 2195 2300 2215
rect 2320 2195 2340 2215
rect 2360 2195 2380 2215
rect 2400 2195 2420 2215
rect 2440 2195 2460 2215
rect 2480 2195 2500 2215
rect 2520 2195 2540 2215
rect 2560 2195 2580 2215
rect 2600 2195 2620 2215
rect 2640 2195 2660 2215
rect 200 2113 220 2133
rect 240 2113 260 2133
rect 280 2113 300 2133
rect 320 2113 340 2133
rect 360 2113 380 2133
rect 400 2113 420 2133
rect 440 2113 460 2133
rect 480 2113 500 2133
rect 520 2113 540 2133
rect 560 2113 580 2133
rect 600 2113 620 2133
rect 640 2113 660 2133
rect 680 2113 700 2133
rect 720 2113 740 2133
rect 760 2113 780 2133
rect 800 2113 820 2133
rect 840 2113 860 2133
rect 880 2113 900 2133
rect 920 2113 940 2133
rect 960 2113 980 2133
rect 1000 2113 1020 2133
rect 1040 2113 1060 2133
rect 1080 2113 1100 2133
rect 1120 2113 1140 2133
rect 1160 2113 1180 2133
rect 1200 2113 1220 2133
rect 1240 2113 1260 2133
rect 1280 2113 1300 2133
rect 1320 2113 1340 2133
rect 1360 2113 1380 2133
rect 1400 2113 1420 2133
rect 1440 2113 1460 2133
rect 1480 2113 1500 2133
rect 1520 2113 1540 2133
rect 1560 2113 1580 2133
rect 1600 2113 1620 2133
rect 1640 2113 1660 2133
rect 1680 2113 1700 2133
rect 1720 2113 1740 2133
rect 1760 2113 1780 2133
rect 1800 2113 1820 2133
rect 1840 2113 1860 2133
rect 1880 2113 1900 2133
rect 1920 2113 1940 2133
rect 1960 2113 1980 2133
rect 2000 2113 2020 2133
rect 2040 2113 2060 2133
rect 2080 2113 2100 2133
rect 2120 2113 2140 2133
rect 2160 2113 2180 2133
rect 2200 2113 2220 2133
rect 2240 2113 2260 2133
rect 2280 2113 2300 2133
rect 2320 2113 2340 2133
rect 2360 2113 2380 2133
rect 2400 2113 2420 2133
rect 2440 2113 2460 2133
rect 2480 2113 2500 2133
rect 2520 2113 2540 2133
rect 2560 2113 2580 2133
rect 2600 2113 2620 2133
rect 2640 2113 2660 2133
rect 200 2031 220 2051
rect 240 2031 260 2051
rect 280 2031 300 2051
rect 320 2031 340 2051
rect 360 2031 380 2051
rect 400 2031 420 2051
rect 440 2031 460 2051
rect 480 2031 500 2051
rect 520 2031 540 2051
rect 560 2031 580 2051
rect 600 2031 620 2051
rect 640 2031 660 2051
rect 680 2031 700 2051
rect 720 2031 740 2051
rect 760 2031 780 2051
rect 800 2031 820 2051
rect 840 2031 860 2051
rect 880 2031 900 2051
rect 920 2031 940 2051
rect 960 2031 980 2051
rect 1000 2031 1020 2051
rect 1040 2031 1060 2051
rect 1080 2031 1100 2051
rect 1120 2031 1140 2051
rect 1160 2031 1180 2051
rect 1200 2031 1220 2051
rect 1240 2031 1260 2051
rect 1280 2031 1300 2051
rect 1320 2031 1340 2051
rect 1360 2031 1380 2051
rect 1400 2031 1420 2051
rect 1440 2031 1460 2051
rect 1480 2031 1500 2051
rect 1520 2031 1540 2051
rect 1560 2031 1580 2051
rect 1600 2031 1620 2051
rect 1640 2031 1660 2051
rect 1680 2031 1700 2051
rect 1720 2031 1740 2051
rect 1760 2031 1780 2051
rect 1800 2031 1820 2051
rect 1840 2031 1860 2051
rect 1880 2031 1900 2051
rect 1920 2031 1940 2051
rect 1960 2031 1980 2051
rect 2000 2031 2020 2051
rect 2040 2031 2060 2051
rect 2080 2031 2100 2051
rect 2120 2031 2140 2051
rect 2160 2031 2180 2051
rect 2200 2031 2220 2051
rect 2240 2031 2260 2051
rect 2280 2031 2300 2051
rect 2320 2031 2340 2051
rect 2360 2031 2380 2051
rect 2400 2031 2420 2051
rect 2440 2031 2460 2051
rect 2480 2031 2500 2051
rect 2520 2031 2540 2051
rect 2560 2031 2580 2051
rect 2600 2031 2620 2051
rect 2640 2031 2660 2051
rect 200 1949 220 1969
rect 240 1949 260 1969
rect 280 1949 300 1969
rect 320 1949 340 1969
rect 360 1949 380 1969
rect 400 1949 420 1969
rect 440 1949 460 1969
rect 480 1949 500 1969
rect 520 1949 540 1969
rect 560 1949 580 1969
rect 600 1949 620 1969
rect 640 1949 660 1969
rect 680 1949 700 1969
rect 720 1949 740 1969
rect 760 1949 780 1969
rect 800 1949 820 1969
rect 840 1949 860 1969
rect 880 1949 900 1969
rect 920 1949 940 1969
rect 960 1949 980 1969
rect 1000 1949 1020 1969
rect 1040 1949 1060 1969
rect 1080 1949 1100 1969
rect 1120 1949 1140 1969
rect 1160 1949 1180 1969
rect 1200 1949 1220 1969
rect 1240 1949 1260 1969
rect 1280 1949 1300 1969
rect 1320 1949 1340 1969
rect 1360 1949 1380 1969
rect 1400 1949 1420 1969
rect 1440 1949 1460 1969
rect 1480 1949 1500 1969
rect 1520 1949 1540 1969
rect 1560 1949 1580 1969
rect 1600 1949 1620 1969
rect 1640 1949 1660 1969
rect 1680 1949 1700 1969
rect 1720 1949 1740 1969
rect 1760 1949 1780 1969
rect 1800 1949 1820 1969
rect 1840 1949 1860 1969
rect 1880 1949 1900 1969
rect 1920 1949 1940 1969
rect 1960 1949 1980 1969
rect 2000 1949 2020 1969
rect 2040 1949 2060 1969
rect 2080 1949 2100 1969
rect 2120 1949 2140 1969
rect 2160 1949 2180 1969
rect 2200 1949 2220 1969
rect 2240 1949 2260 1969
rect 2280 1949 2300 1969
rect 2320 1949 2340 1969
rect 2360 1949 2380 1969
rect 2400 1949 2420 1969
rect 2440 1949 2460 1969
rect 2480 1949 2500 1969
rect 2520 1949 2540 1969
rect 2560 1949 2580 1969
rect 2600 1949 2620 1969
rect 2640 1949 2660 1969
rect 200 1867 220 1887
rect 240 1867 260 1887
rect 280 1867 300 1887
rect 320 1867 340 1887
rect 360 1867 380 1887
rect 400 1867 420 1887
rect 440 1867 460 1887
rect 480 1867 500 1887
rect 520 1867 540 1887
rect 560 1867 580 1887
rect 600 1867 620 1887
rect 640 1867 660 1887
rect 680 1867 700 1887
rect 720 1867 740 1887
rect 760 1867 780 1887
rect 800 1867 820 1887
rect 840 1867 860 1887
rect 880 1867 900 1887
rect 920 1867 940 1887
rect 960 1867 980 1887
rect 1000 1867 1020 1887
rect 1040 1867 1060 1887
rect 1080 1867 1100 1887
rect 1120 1867 1140 1887
rect 1160 1867 1180 1887
rect 1200 1867 1220 1887
rect 1240 1867 1260 1887
rect 1280 1867 1300 1887
rect 1320 1867 1340 1887
rect 1360 1867 1380 1887
rect 1400 1867 1420 1887
rect 1440 1867 1460 1887
rect 1480 1867 1500 1887
rect 1520 1867 1540 1887
rect 1560 1867 1580 1887
rect 1600 1867 1620 1887
rect 1640 1867 1660 1887
rect 1680 1867 1700 1887
rect 1720 1867 1740 1887
rect 1760 1867 1780 1887
rect 1800 1867 1820 1887
rect 1840 1867 1860 1887
rect 1880 1867 1900 1887
rect 1920 1867 1940 1887
rect 1960 1867 1980 1887
rect 2000 1867 2020 1887
rect 2040 1867 2060 1887
rect 2080 1867 2100 1887
rect 2120 1867 2140 1887
rect 2160 1867 2180 1887
rect 2200 1867 2220 1887
rect 2240 1867 2260 1887
rect 2280 1867 2300 1887
rect 2320 1867 2340 1887
rect 2360 1867 2380 1887
rect 2400 1867 2420 1887
rect 2440 1867 2460 1887
rect 2480 1867 2500 1887
rect 2520 1867 2540 1887
rect 2560 1867 2580 1887
rect 2600 1867 2620 1887
rect 2640 1867 2660 1887
rect 200 1785 220 1805
rect 240 1785 260 1805
rect 280 1785 300 1805
rect 320 1785 340 1805
rect 360 1785 380 1805
rect 400 1785 420 1805
rect 440 1785 460 1805
rect 480 1785 500 1805
rect 520 1785 540 1805
rect 560 1785 580 1805
rect 600 1785 620 1805
rect 640 1785 660 1805
rect 680 1785 700 1805
rect 720 1785 740 1805
rect 760 1785 780 1805
rect 800 1785 820 1805
rect 840 1785 860 1805
rect 880 1785 900 1805
rect 920 1785 940 1805
rect 960 1785 980 1805
rect 1000 1785 1020 1805
rect 1040 1785 1060 1805
rect 1080 1785 1100 1805
rect 1120 1785 1140 1805
rect 1160 1785 1180 1805
rect 1200 1785 1220 1805
rect 1240 1785 1260 1805
rect 1280 1785 1300 1805
rect 1320 1785 1340 1805
rect 1360 1785 1380 1805
rect 1400 1785 1420 1805
rect 1440 1785 1460 1805
rect 1480 1785 1500 1805
rect 1520 1785 1540 1805
rect 1560 1785 1580 1805
rect 1600 1785 1620 1805
rect 1640 1785 1660 1805
rect 1680 1785 1700 1805
rect 1720 1785 1740 1805
rect 1760 1785 1780 1805
rect 1800 1785 1820 1805
rect 1840 1785 1860 1805
rect 1880 1785 1900 1805
rect 1920 1785 1940 1805
rect 1960 1785 1980 1805
rect 2000 1785 2020 1805
rect 2040 1785 2060 1805
rect 2080 1785 2100 1805
rect 2120 1785 2140 1805
rect 2160 1785 2180 1805
rect 2200 1785 2220 1805
rect 2240 1785 2260 1805
rect 2280 1785 2300 1805
rect 2320 1785 2340 1805
rect 2360 1785 2380 1805
rect 2400 1785 2420 1805
rect 2440 1785 2460 1805
rect 2480 1785 2500 1805
rect 2520 1785 2540 1805
rect 2560 1785 2580 1805
rect 2600 1785 2620 1805
rect 2640 1785 2660 1805
rect 200 1703 220 1723
rect 240 1703 260 1723
rect 280 1703 300 1723
rect 320 1703 340 1723
rect 360 1703 380 1723
rect 400 1703 420 1723
rect 440 1703 460 1723
rect 480 1703 500 1723
rect 520 1703 540 1723
rect 560 1703 580 1723
rect 600 1703 620 1723
rect 640 1703 660 1723
rect 680 1703 700 1723
rect 720 1703 740 1723
rect 760 1703 780 1723
rect 800 1703 820 1723
rect 840 1703 860 1723
rect 880 1703 900 1723
rect 920 1703 940 1723
rect 960 1703 980 1723
rect 1000 1703 1020 1723
rect 1040 1703 1060 1723
rect 1080 1703 1100 1723
rect 1120 1703 1140 1723
rect 1160 1703 1180 1723
rect 1200 1703 1220 1723
rect 1240 1703 1260 1723
rect 1280 1703 1300 1723
rect 1320 1703 1340 1723
rect 1360 1703 1380 1723
rect 1400 1703 1420 1723
rect 1440 1703 1460 1723
rect 1480 1703 1500 1723
rect 1520 1703 1540 1723
rect 1560 1703 1580 1723
rect 1600 1703 1620 1723
rect 1640 1703 1660 1723
rect 1680 1703 1700 1723
rect 1720 1703 1740 1723
rect 1760 1703 1780 1723
rect 1800 1703 1820 1723
rect 1840 1703 1860 1723
rect 1880 1703 1900 1723
rect 1920 1703 1940 1723
rect 1960 1703 1980 1723
rect 2000 1703 2020 1723
rect 2040 1703 2060 1723
rect 2080 1703 2100 1723
rect 2120 1703 2140 1723
rect 2160 1703 2180 1723
rect 2200 1703 2220 1723
rect 2240 1703 2260 1723
rect 2280 1703 2300 1723
rect 2320 1703 2340 1723
rect 2360 1703 2380 1723
rect 2400 1703 2420 1723
rect 2440 1703 2460 1723
rect 2480 1703 2500 1723
rect 2520 1703 2540 1723
rect 2560 1703 2580 1723
rect 2600 1703 2620 1723
rect 2640 1703 2660 1723
rect 200 1621 220 1641
rect 240 1621 260 1641
rect 280 1621 300 1641
rect 320 1621 340 1641
rect 360 1621 380 1641
rect 400 1621 420 1641
rect 440 1621 460 1641
rect 480 1621 500 1641
rect 520 1621 540 1641
rect 560 1621 580 1641
rect 600 1621 620 1641
rect 640 1621 660 1641
rect 680 1621 700 1641
rect 720 1621 740 1641
rect 760 1621 780 1641
rect 800 1621 820 1641
rect 840 1621 860 1641
rect 880 1621 900 1641
rect 920 1621 940 1641
rect 960 1621 980 1641
rect 1000 1621 1020 1641
rect 1040 1621 1060 1641
rect 1080 1621 1100 1641
rect 1120 1621 1140 1641
rect 1160 1621 1180 1641
rect 1200 1621 1220 1641
rect 1240 1621 1260 1641
rect 1280 1621 1300 1641
rect 1320 1621 1340 1641
rect 1360 1621 1380 1641
rect 1400 1621 1420 1641
rect 1440 1621 1460 1641
rect 1480 1621 1500 1641
rect 1520 1621 1540 1641
rect 1560 1621 1580 1641
rect 1600 1621 1620 1641
rect 1640 1621 1660 1641
rect 1680 1621 1700 1641
rect 1720 1621 1740 1641
rect 1760 1621 1780 1641
rect 1800 1621 1820 1641
rect 1840 1621 1860 1641
rect 1880 1621 1900 1641
rect 1920 1621 1940 1641
rect 1960 1621 1980 1641
rect 2000 1621 2020 1641
rect 2040 1621 2060 1641
rect 2080 1621 2100 1641
rect 2120 1621 2140 1641
rect 2160 1621 2180 1641
rect 2200 1621 2220 1641
rect 2240 1621 2260 1641
rect 2280 1621 2300 1641
rect 2320 1621 2340 1641
rect 2360 1621 2380 1641
rect 2400 1621 2420 1641
rect 2440 1621 2460 1641
rect 2480 1621 2500 1641
rect 2520 1621 2540 1641
rect 2560 1621 2580 1641
rect 2600 1621 2620 1641
rect 2640 1621 2660 1641
rect 200 1539 220 1559
rect 240 1539 260 1559
rect 280 1539 300 1559
rect 320 1539 340 1559
rect 360 1539 380 1559
rect 400 1539 420 1559
rect 440 1539 460 1559
rect 480 1539 500 1559
rect 520 1539 540 1559
rect 560 1539 580 1559
rect 600 1539 620 1559
rect 640 1539 660 1559
rect 680 1539 700 1559
rect 720 1539 740 1559
rect 760 1539 780 1559
rect 800 1539 820 1559
rect 840 1539 860 1559
rect 880 1539 900 1559
rect 920 1539 940 1559
rect 960 1539 980 1559
rect 1000 1539 1020 1559
rect 1040 1539 1060 1559
rect 1080 1539 1100 1559
rect 1120 1539 1140 1559
rect 1160 1539 1180 1559
rect 1200 1539 1220 1559
rect 1240 1539 1260 1559
rect 1280 1539 1300 1559
rect 1320 1539 1340 1559
rect 1360 1539 1380 1559
rect 1400 1539 1420 1559
rect 1440 1539 1460 1559
rect 1480 1539 1500 1559
rect 1520 1539 1540 1559
rect 1560 1539 1580 1559
rect 1600 1539 1620 1559
rect 1640 1539 1660 1559
rect 1680 1539 1700 1559
rect 1720 1539 1740 1559
rect 1760 1539 1780 1559
rect 1800 1539 1820 1559
rect 1840 1539 1860 1559
rect 1880 1539 1900 1559
rect 1920 1539 1940 1559
rect 1960 1539 1980 1559
rect 2000 1539 2020 1559
rect 2040 1539 2060 1559
rect 2080 1539 2100 1559
rect 2120 1539 2140 1559
rect 2160 1539 2180 1559
rect 2200 1539 2220 1559
rect 2240 1539 2260 1559
rect 2280 1539 2300 1559
rect 2320 1539 2340 1559
rect 2360 1539 2380 1559
rect 2400 1539 2420 1559
rect 2440 1539 2460 1559
rect 2480 1539 2500 1559
rect 2520 1539 2540 1559
rect 2560 1539 2580 1559
rect 2600 1539 2620 1559
rect 2640 1539 2660 1559
rect 200 1457 220 1477
rect 240 1457 260 1477
rect 280 1457 300 1477
rect 320 1457 340 1477
rect 360 1457 380 1477
rect 400 1457 420 1477
rect 440 1457 460 1477
rect 480 1457 500 1477
rect 520 1457 540 1477
rect 560 1457 580 1477
rect 600 1457 620 1477
rect 640 1457 660 1477
rect 680 1457 700 1477
rect 720 1457 740 1477
rect 760 1457 780 1477
rect 800 1457 820 1477
rect 840 1457 860 1477
rect 880 1457 900 1477
rect 920 1457 940 1477
rect 960 1457 980 1477
rect 1000 1457 1020 1477
rect 1040 1457 1060 1477
rect 1080 1457 1100 1477
rect 1120 1457 1140 1477
rect 1160 1457 1180 1477
rect 1200 1457 1220 1477
rect 1240 1457 1260 1477
rect 1280 1457 1300 1477
rect 1320 1457 1340 1477
rect 1360 1457 1380 1477
rect 1400 1457 1420 1477
rect 1440 1457 1460 1477
rect 1480 1457 1500 1477
rect 1520 1457 1540 1477
rect 1560 1457 1580 1477
rect 1600 1457 1620 1477
rect 1640 1457 1660 1477
rect 1680 1457 1700 1477
rect 1720 1457 1740 1477
rect 1760 1457 1780 1477
rect 1800 1457 1820 1477
rect 1840 1457 1860 1477
rect 1880 1457 1900 1477
rect 1920 1457 1940 1477
rect 1960 1457 1980 1477
rect 2000 1457 2020 1477
rect 2040 1457 2060 1477
rect 2080 1457 2100 1477
rect 2120 1457 2140 1477
rect 2160 1457 2180 1477
rect 2200 1457 2220 1477
rect 2240 1457 2260 1477
rect 2280 1457 2300 1477
rect 2320 1457 2340 1477
rect 2360 1457 2380 1477
rect 2400 1457 2420 1477
rect 2440 1457 2460 1477
rect 2480 1457 2500 1477
rect 2520 1457 2540 1477
rect 2560 1457 2580 1477
rect 2600 1457 2620 1477
rect 2640 1457 2660 1477
rect 200 1375 220 1395
rect 240 1375 260 1395
rect 280 1375 300 1395
rect 320 1375 340 1395
rect 360 1375 380 1395
rect 400 1375 420 1395
rect 440 1375 460 1395
rect 480 1375 500 1395
rect 520 1375 540 1395
rect 560 1375 580 1395
rect 600 1375 620 1395
rect 640 1375 660 1395
rect 680 1375 700 1395
rect 720 1375 740 1395
rect 760 1375 780 1395
rect 800 1375 820 1395
rect 840 1375 860 1395
rect 880 1375 900 1395
rect 920 1375 940 1395
rect 960 1375 980 1395
rect 1000 1375 1020 1395
rect 1040 1375 1060 1395
rect 1080 1375 1100 1395
rect 1120 1375 1140 1395
rect 1160 1375 1180 1395
rect 1200 1375 1220 1395
rect 1240 1375 1260 1395
rect 1280 1375 1300 1395
rect 1320 1375 1340 1395
rect 1360 1375 1380 1395
rect 1400 1375 1420 1395
rect 1440 1375 1460 1395
rect 1480 1375 1500 1395
rect 1520 1375 1540 1395
rect 1560 1375 1580 1395
rect 1600 1375 1620 1395
rect 1640 1375 1660 1395
rect 1680 1375 1700 1395
rect 1720 1375 1740 1395
rect 1760 1375 1780 1395
rect 1800 1375 1820 1395
rect 1840 1375 1860 1395
rect 1880 1375 1900 1395
rect 1920 1375 1940 1395
rect 1960 1375 1980 1395
rect 2000 1375 2020 1395
rect 2040 1375 2060 1395
rect 2080 1375 2100 1395
rect 2120 1375 2140 1395
rect 2160 1375 2180 1395
rect 2200 1375 2220 1395
rect 2240 1375 2260 1395
rect 2280 1375 2300 1395
rect 2320 1375 2340 1395
rect 2360 1375 2380 1395
rect 2400 1375 2420 1395
rect 2440 1375 2460 1395
rect 2480 1375 2500 1395
rect 2520 1375 2540 1395
rect 2560 1375 2580 1395
rect 2600 1375 2620 1395
rect 2640 1375 2660 1395
rect 200 1293 220 1313
rect 240 1293 260 1313
rect 280 1293 300 1313
rect 320 1293 340 1313
rect 360 1293 380 1313
rect 400 1293 420 1313
rect 440 1293 460 1313
rect 480 1293 500 1313
rect 520 1293 540 1313
rect 560 1293 580 1313
rect 600 1293 620 1313
rect 640 1293 660 1313
rect 680 1293 700 1313
rect 720 1293 740 1313
rect 760 1293 780 1313
rect 800 1293 820 1313
rect 840 1293 860 1313
rect 880 1293 900 1313
rect 920 1293 940 1313
rect 960 1293 980 1313
rect 1000 1293 1020 1313
rect 1040 1293 1060 1313
rect 1080 1293 1100 1313
rect 1120 1293 1140 1313
rect 1160 1293 1180 1313
rect 1200 1293 1220 1313
rect 1240 1293 1260 1313
rect 1280 1293 1300 1313
rect 1320 1293 1340 1313
rect 1360 1293 1380 1313
rect 1400 1293 1420 1313
rect 1440 1293 1460 1313
rect 1480 1293 1500 1313
rect 1520 1293 1540 1313
rect 1560 1293 1580 1313
rect 1600 1293 1620 1313
rect 1640 1293 1660 1313
rect 1680 1293 1700 1313
rect 1720 1293 1740 1313
rect 1760 1293 1780 1313
rect 1800 1293 1820 1313
rect 1840 1293 1860 1313
rect 1880 1293 1900 1313
rect 1920 1293 1940 1313
rect 1960 1293 1980 1313
rect 2000 1293 2020 1313
rect 2040 1293 2060 1313
rect 2080 1293 2100 1313
rect 2120 1293 2140 1313
rect 2160 1293 2180 1313
rect 2200 1293 2220 1313
rect 2240 1293 2260 1313
rect 2280 1293 2300 1313
rect 2320 1293 2340 1313
rect 2360 1293 2380 1313
rect 2400 1293 2420 1313
rect 2440 1293 2460 1313
rect 2480 1293 2500 1313
rect 2520 1293 2540 1313
rect 2560 1293 2580 1313
rect 2600 1293 2620 1313
rect 2640 1293 2660 1313
rect 200 1211 220 1231
rect 240 1211 260 1231
rect 280 1211 300 1231
rect 320 1211 340 1231
rect 360 1211 380 1231
rect 400 1211 420 1231
rect 440 1211 460 1231
rect 480 1211 500 1231
rect 520 1211 540 1231
rect 560 1211 580 1231
rect 600 1211 620 1231
rect 640 1211 660 1231
rect 680 1211 700 1231
rect 720 1211 740 1231
rect 760 1211 780 1231
rect 800 1211 820 1231
rect 840 1211 860 1231
rect 880 1211 900 1231
rect 920 1211 940 1231
rect 960 1211 980 1231
rect 1000 1211 1020 1231
rect 1040 1211 1060 1231
rect 1080 1211 1100 1231
rect 1120 1211 1140 1231
rect 1160 1211 1180 1231
rect 1200 1211 1220 1231
rect 1240 1211 1260 1231
rect 1280 1211 1300 1231
rect 1320 1211 1340 1231
rect 1360 1211 1380 1231
rect 1400 1211 1420 1231
rect 1440 1211 1460 1231
rect 1480 1211 1500 1231
rect 1520 1211 1540 1231
rect 1560 1211 1580 1231
rect 1600 1211 1620 1231
rect 1640 1211 1660 1231
rect 1680 1211 1700 1231
rect 1720 1211 1740 1231
rect 1760 1211 1780 1231
rect 1800 1211 1820 1231
rect 1840 1211 1860 1231
rect 1880 1211 1900 1231
rect 1920 1211 1940 1231
rect 1960 1211 1980 1231
rect 2000 1211 2020 1231
rect 2040 1211 2060 1231
rect 2080 1211 2100 1231
rect 2120 1211 2140 1231
rect 2160 1211 2180 1231
rect 2200 1211 2220 1231
rect 2240 1211 2260 1231
rect 2280 1211 2300 1231
rect 2320 1211 2340 1231
rect 2360 1211 2380 1231
rect 2400 1211 2420 1231
rect 2440 1211 2460 1231
rect 2480 1211 2500 1231
rect 2520 1211 2540 1231
rect 2560 1211 2580 1231
rect 2600 1211 2620 1231
rect 2640 1211 2660 1231
rect 200 1129 220 1149
rect 240 1129 260 1149
rect 280 1129 300 1149
rect 320 1129 340 1149
rect 360 1129 380 1149
rect 400 1129 420 1149
rect 440 1129 460 1149
rect 480 1129 500 1149
rect 520 1129 540 1149
rect 560 1129 580 1149
rect 600 1129 620 1149
rect 640 1129 660 1149
rect 680 1129 700 1149
rect 720 1129 740 1149
rect 760 1129 780 1149
rect 800 1129 820 1149
rect 840 1129 860 1149
rect 880 1129 900 1149
rect 920 1129 940 1149
rect 960 1129 980 1149
rect 1000 1129 1020 1149
rect 1040 1129 1060 1149
rect 1080 1129 1100 1149
rect 1120 1129 1140 1149
rect 1160 1129 1180 1149
rect 1200 1129 1220 1149
rect 1240 1129 1260 1149
rect 1280 1129 1300 1149
rect 1320 1129 1340 1149
rect 1360 1129 1380 1149
rect 1400 1129 1420 1149
rect 1440 1129 1460 1149
rect 1480 1129 1500 1149
rect 1520 1129 1540 1149
rect 1560 1129 1580 1149
rect 1600 1129 1620 1149
rect 1640 1129 1660 1149
rect 1680 1129 1700 1149
rect 1720 1129 1740 1149
rect 1760 1129 1780 1149
rect 1800 1129 1820 1149
rect 1840 1129 1860 1149
rect 1880 1129 1900 1149
rect 1920 1129 1940 1149
rect 1960 1129 1980 1149
rect 2000 1129 2020 1149
rect 2040 1129 2060 1149
rect 2080 1129 2100 1149
rect 2120 1129 2140 1149
rect 2160 1129 2180 1149
rect 2200 1129 2220 1149
rect 2240 1129 2260 1149
rect 2280 1129 2300 1149
rect 2320 1129 2340 1149
rect 2360 1129 2380 1149
rect 2400 1129 2420 1149
rect 2440 1129 2460 1149
rect 2480 1129 2500 1149
rect 2520 1129 2540 1149
rect 2560 1129 2580 1149
rect 2600 1129 2620 1149
rect 2640 1129 2660 1149
rect 200 1047 220 1067
rect 240 1047 260 1067
rect 280 1047 300 1067
rect 320 1047 340 1067
rect 360 1047 380 1067
rect 400 1047 420 1067
rect 440 1047 460 1067
rect 480 1047 500 1067
rect 520 1047 540 1067
rect 560 1047 580 1067
rect 600 1047 620 1067
rect 640 1047 660 1067
rect 680 1047 700 1067
rect 720 1047 740 1067
rect 760 1047 780 1067
rect 800 1047 820 1067
rect 840 1047 860 1067
rect 880 1047 900 1067
rect 920 1047 940 1067
rect 960 1047 980 1067
rect 1000 1047 1020 1067
rect 1040 1047 1060 1067
rect 1080 1047 1100 1067
rect 1120 1047 1140 1067
rect 1160 1047 1180 1067
rect 1200 1047 1220 1067
rect 1240 1047 1260 1067
rect 1280 1047 1300 1067
rect 1320 1047 1340 1067
rect 1360 1047 1380 1067
rect 1400 1047 1420 1067
rect 1440 1047 1460 1067
rect 1480 1047 1500 1067
rect 1520 1047 1540 1067
rect 1560 1047 1580 1067
rect 1600 1047 1620 1067
rect 1640 1047 1660 1067
rect 1680 1047 1700 1067
rect 1720 1047 1740 1067
rect 1760 1047 1780 1067
rect 1800 1047 1820 1067
rect 1840 1047 1860 1067
rect 1880 1047 1900 1067
rect 1920 1047 1940 1067
rect 1960 1047 1980 1067
rect 2000 1047 2020 1067
rect 2040 1047 2060 1067
rect 2080 1047 2100 1067
rect 2120 1047 2140 1067
rect 2160 1047 2180 1067
rect 2200 1047 2220 1067
rect 2240 1047 2260 1067
rect 2280 1047 2300 1067
rect 2320 1047 2340 1067
rect 2360 1047 2380 1067
rect 2400 1047 2420 1067
rect 2440 1047 2460 1067
rect 2480 1047 2500 1067
rect 2520 1047 2540 1067
rect 2560 1047 2580 1067
rect 2600 1047 2620 1067
rect 2640 1047 2660 1067
rect 200 965 220 985
rect 240 965 260 985
rect 280 965 300 985
rect 320 965 340 985
rect 360 965 380 985
rect 400 965 420 985
rect 440 965 460 985
rect 480 965 500 985
rect 520 965 540 985
rect 560 965 580 985
rect 600 965 620 985
rect 640 965 660 985
rect 680 965 700 985
rect 720 965 740 985
rect 760 965 780 985
rect 800 965 820 985
rect 840 965 860 985
rect 880 965 900 985
rect 920 965 940 985
rect 960 965 980 985
rect 1000 965 1020 985
rect 1040 965 1060 985
rect 1080 965 1100 985
rect 1120 965 1140 985
rect 1160 965 1180 985
rect 1200 965 1220 985
rect 1240 965 1260 985
rect 1280 965 1300 985
rect 1320 965 1340 985
rect 1360 965 1380 985
rect 1400 965 1420 985
rect 1440 965 1460 985
rect 1480 965 1500 985
rect 1520 965 1540 985
rect 1560 965 1580 985
rect 1600 965 1620 985
rect 1640 965 1660 985
rect 1680 965 1700 985
rect 1720 965 1740 985
rect 1760 965 1780 985
rect 1800 965 1820 985
rect 1840 965 1860 985
rect 1880 965 1900 985
rect 1920 965 1940 985
rect 1960 965 1980 985
rect 2000 965 2020 985
rect 2040 965 2060 985
rect 2080 965 2100 985
rect 2120 965 2140 985
rect 2160 965 2180 985
rect 2200 965 2220 985
rect 2240 965 2260 985
rect 2280 965 2300 985
rect 2320 965 2340 985
rect 2360 965 2380 985
rect 2400 965 2420 985
rect 2440 965 2460 985
rect 2480 965 2500 985
rect 2520 965 2540 985
rect 2560 965 2580 985
rect 2600 965 2620 985
rect 2640 965 2660 985
rect 200 883 220 903
rect 240 883 260 903
rect 280 883 300 903
rect 320 883 340 903
rect 360 883 380 903
rect 400 883 420 903
rect 440 883 460 903
rect 480 883 500 903
rect 520 883 540 903
rect 560 883 580 903
rect 600 883 620 903
rect 640 883 660 903
rect 680 883 700 903
rect 720 883 740 903
rect 760 883 780 903
rect 800 883 820 903
rect 840 883 860 903
rect 880 883 900 903
rect 920 883 940 903
rect 960 883 980 903
rect 1000 883 1020 903
rect 1040 883 1060 903
rect 1080 883 1100 903
rect 1120 883 1140 903
rect 1160 883 1180 903
rect 1200 883 1220 903
rect 1240 883 1260 903
rect 1280 883 1300 903
rect 1320 883 1340 903
rect 1360 883 1380 903
rect 1400 883 1420 903
rect 1440 883 1460 903
rect 1480 883 1500 903
rect 1520 883 1540 903
rect 1560 883 1580 903
rect 1600 883 1620 903
rect 1640 883 1660 903
rect 1680 883 1700 903
rect 1720 883 1740 903
rect 1760 883 1780 903
rect 1800 883 1820 903
rect 1840 883 1860 903
rect 1880 883 1900 903
rect 1920 883 1940 903
rect 1960 883 1980 903
rect 2000 883 2020 903
rect 2040 883 2060 903
rect 2080 883 2100 903
rect 2120 883 2140 903
rect 2160 883 2180 903
rect 2200 883 2220 903
rect 2240 883 2260 903
rect 2280 883 2300 903
rect 2320 883 2340 903
rect 2360 883 2380 903
rect 2400 883 2420 903
rect 2440 883 2460 903
rect 2480 883 2500 903
rect 2520 883 2540 903
rect 2560 883 2580 903
rect 2600 883 2620 903
rect 2640 883 2660 903
rect 200 801 220 821
rect 240 801 260 821
rect 280 801 300 821
rect 320 801 340 821
rect 360 801 380 821
rect 400 801 420 821
rect 440 801 460 821
rect 480 801 500 821
rect 520 801 540 821
rect 560 801 580 821
rect 600 801 620 821
rect 640 801 660 821
rect 680 801 700 821
rect 720 801 740 821
rect 760 801 780 821
rect 800 801 820 821
rect 840 801 860 821
rect 880 801 900 821
rect 920 801 940 821
rect 960 801 980 821
rect 1000 801 1020 821
rect 1040 801 1060 821
rect 1080 801 1100 821
rect 1120 801 1140 821
rect 1160 801 1180 821
rect 1200 801 1220 821
rect 1240 801 1260 821
rect 1280 801 1300 821
rect 1320 801 1340 821
rect 1360 801 1380 821
rect 1400 801 1420 821
rect 1440 801 1460 821
rect 1480 801 1500 821
rect 1520 801 1540 821
rect 1560 801 1580 821
rect 1600 801 1620 821
rect 1640 801 1660 821
rect 1680 801 1700 821
rect 1720 801 1740 821
rect 1760 801 1780 821
rect 1800 801 1820 821
rect 1840 801 1860 821
rect 1880 801 1900 821
rect 1920 801 1940 821
rect 1960 801 1980 821
rect 2000 801 2020 821
rect 2040 801 2060 821
rect 2080 801 2100 821
rect 2120 801 2140 821
rect 2160 801 2180 821
rect 2200 801 2220 821
rect 2240 801 2260 821
rect 2280 801 2300 821
rect 2320 801 2340 821
rect 2360 801 2380 821
rect 2400 801 2420 821
rect 2440 801 2460 821
rect 2480 801 2500 821
rect 2520 801 2540 821
rect 2560 801 2580 821
rect 2600 801 2620 821
rect 2640 801 2660 821
rect 200 719 220 739
rect 240 719 260 739
rect 280 719 300 739
rect 320 719 340 739
rect 360 719 380 739
rect 400 719 420 739
rect 440 719 460 739
rect 480 719 500 739
rect 520 719 540 739
rect 560 719 580 739
rect 600 719 620 739
rect 640 719 660 739
rect 680 719 700 739
rect 720 719 740 739
rect 760 719 780 739
rect 800 719 820 739
rect 840 719 860 739
rect 880 719 900 739
rect 920 719 940 739
rect 960 719 980 739
rect 1000 719 1020 739
rect 1040 719 1060 739
rect 1080 719 1100 739
rect 1120 719 1140 739
rect 1160 719 1180 739
rect 1200 719 1220 739
rect 1240 719 1260 739
rect 1280 719 1300 739
rect 1320 719 1340 739
rect 1360 719 1380 739
rect 1400 719 1420 739
rect 1440 719 1460 739
rect 1480 719 1500 739
rect 1520 719 1540 739
rect 1560 719 1580 739
rect 1600 719 1620 739
rect 1640 719 1660 739
rect 1680 719 1700 739
rect 1720 719 1740 739
rect 1760 719 1780 739
rect 1800 719 1820 739
rect 1840 719 1860 739
rect 1880 719 1900 739
rect 1920 719 1940 739
rect 1960 719 1980 739
rect 2000 719 2020 739
rect 2040 719 2060 739
rect 2080 719 2100 739
rect 2120 719 2140 739
rect 2160 719 2180 739
rect 2200 719 2220 739
rect 2240 719 2260 739
rect 2280 719 2300 739
rect 2320 719 2340 739
rect 2360 719 2380 739
rect 2400 719 2420 739
rect 2440 719 2460 739
rect 2480 719 2500 739
rect 2520 719 2540 739
rect 2560 719 2580 739
rect 2600 719 2620 739
rect 2640 719 2660 739
rect 200 637 220 657
rect 240 637 260 657
rect 280 637 300 657
rect 320 637 340 657
rect 360 637 380 657
rect 400 637 420 657
rect 440 637 460 657
rect 480 637 500 657
rect 520 637 540 657
rect 560 637 580 657
rect 600 637 620 657
rect 640 637 660 657
rect 680 637 700 657
rect 720 637 740 657
rect 760 637 780 657
rect 800 637 820 657
rect 840 637 860 657
rect 880 637 900 657
rect 920 637 940 657
rect 960 637 980 657
rect 1000 637 1020 657
rect 1040 637 1060 657
rect 1080 637 1100 657
rect 1120 637 1140 657
rect 1160 637 1180 657
rect 1200 637 1220 657
rect 1240 637 1260 657
rect 1280 637 1300 657
rect 1320 637 1340 657
rect 1360 637 1380 657
rect 1400 637 1420 657
rect 1440 637 1460 657
rect 1480 637 1500 657
rect 1520 637 1540 657
rect 1560 637 1580 657
rect 1600 637 1620 657
rect 1640 637 1660 657
rect 1680 637 1700 657
rect 1720 637 1740 657
rect 1760 637 1780 657
rect 1800 637 1820 657
rect 1840 637 1860 657
rect 1880 637 1900 657
rect 1920 637 1940 657
rect 1960 637 1980 657
rect 2000 637 2020 657
rect 2040 637 2060 657
rect 2080 637 2100 657
rect 2120 637 2140 657
rect 2160 637 2180 657
rect 2200 637 2220 657
rect 2240 637 2260 657
rect 2280 637 2300 657
rect 2320 637 2340 657
rect 2360 637 2380 657
rect 2400 637 2420 657
rect 2440 637 2460 657
rect 2480 637 2500 657
rect 2520 637 2540 657
rect 2560 637 2580 657
rect 2600 637 2620 657
rect 2640 637 2660 657
rect 200 555 220 575
rect 240 555 260 575
rect 280 555 300 575
rect 320 555 340 575
rect 360 555 380 575
rect 400 555 420 575
rect 440 555 460 575
rect 480 555 500 575
rect 520 555 540 575
rect 560 555 580 575
rect 600 555 620 575
rect 640 555 660 575
rect 680 555 700 575
rect 720 555 740 575
rect 760 555 780 575
rect 800 555 820 575
rect 840 555 860 575
rect 880 555 900 575
rect 920 555 940 575
rect 960 555 980 575
rect 1000 555 1020 575
rect 1040 555 1060 575
rect 1080 555 1100 575
rect 1120 555 1140 575
rect 1160 555 1180 575
rect 1200 555 1220 575
rect 1240 555 1260 575
rect 1280 555 1300 575
rect 1320 555 1340 575
rect 1360 555 1380 575
rect 1400 555 1420 575
rect 1440 555 1460 575
rect 1480 555 1500 575
rect 1520 555 1540 575
rect 1560 555 1580 575
rect 1600 555 1620 575
rect 1640 555 1660 575
rect 1680 555 1700 575
rect 1720 555 1740 575
rect 1760 555 1780 575
rect 1800 555 1820 575
rect 1840 555 1860 575
rect 1880 555 1900 575
rect 1920 555 1940 575
rect 1960 555 1980 575
rect 2000 555 2020 575
rect 2040 555 2060 575
rect 2080 555 2100 575
rect 2120 555 2140 575
rect 2160 555 2180 575
rect 2200 555 2220 575
rect 2240 555 2260 575
rect 2280 555 2300 575
rect 2320 555 2340 575
rect 2360 555 2380 575
rect 2400 555 2420 575
rect 2440 555 2460 575
rect 2480 555 2500 575
rect 2520 555 2540 575
rect 2560 555 2580 575
rect 2600 555 2620 575
rect 2640 555 2660 575
rect 200 473 220 493
rect 240 473 260 493
rect 280 473 300 493
rect 320 473 340 493
rect 360 473 380 493
rect 400 473 420 493
rect 440 473 460 493
rect 480 473 500 493
rect 520 473 540 493
rect 560 473 580 493
rect 600 473 620 493
rect 640 473 660 493
rect 680 473 700 493
rect 720 473 740 493
rect 760 473 780 493
rect 800 473 820 493
rect 840 473 860 493
rect 880 473 900 493
rect 920 473 940 493
rect 960 473 980 493
rect 1000 473 1020 493
rect 1040 473 1060 493
rect 1080 473 1100 493
rect 1120 473 1140 493
rect 1160 473 1180 493
rect 1200 473 1220 493
rect 1240 473 1260 493
rect 1280 473 1300 493
rect 1320 473 1340 493
rect 1360 473 1380 493
rect 1400 473 1420 493
rect 1440 473 1460 493
rect 1480 473 1500 493
rect 1520 473 1540 493
rect 1560 473 1580 493
rect 1600 473 1620 493
rect 1640 473 1660 493
rect 1680 473 1700 493
rect 1720 473 1740 493
rect 1760 473 1780 493
rect 1800 473 1820 493
rect 1840 473 1860 493
rect 1880 473 1900 493
rect 1920 473 1940 493
rect 1960 473 1980 493
rect 2000 473 2020 493
rect 2040 473 2060 493
rect 2080 473 2100 493
rect 2120 473 2140 493
rect 2160 473 2180 493
rect 2200 473 2220 493
rect 2240 473 2260 493
rect 2280 473 2300 493
rect 2320 473 2340 493
rect 2360 473 2380 493
rect 2400 473 2420 493
rect 2440 473 2460 493
rect 2480 473 2500 493
rect 2520 473 2540 493
rect 2560 473 2580 493
rect 2600 473 2620 493
rect 2640 473 2660 493
rect 200 391 220 411
rect 240 391 260 411
rect 280 391 300 411
rect 320 391 340 411
rect 360 391 380 411
rect 400 391 420 411
rect 440 391 460 411
rect 480 391 500 411
rect 520 391 540 411
rect 560 391 580 411
rect 600 391 620 411
rect 640 391 660 411
rect 680 391 700 411
rect 720 391 740 411
rect 760 391 780 411
rect 800 391 820 411
rect 840 391 860 411
rect 880 391 900 411
rect 920 391 940 411
rect 960 391 980 411
rect 1000 391 1020 411
rect 1040 391 1060 411
rect 1080 391 1100 411
rect 1120 391 1140 411
rect 1160 391 1180 411
rect 1200 391 1220 411
rect 1240 391 1260 411
rect 1280 391 1300 411
rect 1320 391 1340 411
rect 1360 391 1380 411
rect 1400 391 1420 411
rect 1440 391 1460 411
rect 1480 391 1500 411
rect 1520 391 1540 411
rect 1560 391 1580 411
rect 1600 391 1620 411
rect 1640 391 1660 411
rect 1680 391 1700 411
rect 1720 391 1740 411
rect 1760 391 1780 411
rect 1800 391 1820 411
rect 1840 391 1860 411
rect 1880 391 1900 411
rect 1920 391 1940 411
rect 1960 391 1980 411
rect 2000 391 2020 411
rect 2040 391 2060 411
rect 2080 391 2100 411
rect 2120 391 2140 411
rect 2160 391 2180 411
rect 2200 391 2220 411
rect 2240 391 2260 411
rect 2280 391 2300 411
rect 2320 391 2340 411
rect 2360 391 2380 411
rect 2400 391 2420 411
rect 2440 391 2460 411
rect 2480 391 2500 411
rect 2520 391 2540 411
rect 2560 391 2580 411
rect 2600 391 2620 411
rect 2640 391 2660 411
rect 200 309 220 329
rect 240 309 260 329
rect 280 309 300 329
rect 320 309 340 329
rect 360 309 380 329
rect 400 309 420 329
rect 440 309 460 329
rect 480 309 500 329
rect 520 309 540 329
rect 560 309 580 329
rect 600 309 620 329
rect 640 309 660 329
rect 680 309 700 329
rect 720 309 740 329
rect 760 309 780 329
rect 800 309 820 329
rect 840 309 860 329
rect 880 309 900 329
rect 920 309 940 329
rect 960 309 980 329
rect 1000 309 1020 329
rect 1040 309 1060 329
rect 1080 309 1100 329
rect 1120 309 1140 329
rect 1160 309 1180 329
rect 1200 309 1220 329
rect 1240 309 1260 329
rect 1280 309 1300 329
rect 1320 309 1340 329
rect 1360 309 1380 329
rect 1400 309 1420 329
rect 1440 309 1460 329
rect 1480 309 1500 329
rect 1520 309 1540 329
rect 1560 309 1580 329
rect 1600 309 1620 329
rect 1640 309 1660 329
rect 1680 309 1700 329
rect 1720 309 1740 329
rect 1760 309 1780 329
rect 1800 309 1820 329
rect 1840 309 1860 329
rect 1880 309 1900 329
rect 1920 309 1940 329
rect 1960 309 1980 329
rect 2000 309 2020 329
rect 2040 309 2060 329
rect 2080 309 2100 329
rect 2120 309 2140 329
rect 2160 309 2180 329
rect 2200 309 2220 329
rect 2240 309 2260 329
rect 2280 309 2300 329
rect 2320 309 2340 329
rect 2360 309 2380 329
rect 2400 309 2420 329
rect 2440 309 2460 329
rect 2480 309 2500 329
rect 2520 309 2540 329
rect 2560 309 2580 329
rect 2600 309 2620 329
rect 2640 309 2660 329
rect 200 227 220 247
rect 240 227 260 247
rect 280 227 300 247
rect 320 227 340 247
rect 360 227 380 247
rect 400 227 420 247
rect 440 227 460 247
rect 480 227 500 247
rect 520 227 540 247
rect 560 227 580 247
rect 600 227 620 247
rect 640 227 660 247
rect 680 227 700 247
rect 720 227 740 247
rect 760 227 780 247
rect 800 227 820 247
rect 840 227 860 247
rect 880 227 900 247
rect 920 227 940 247
rect 960 227 980 247
rect 1000 227 1020 247
rect 1040 227 1060 247
rect 1080 227 1100 247
rect 1120 227 1140 247
rect 1160 227 1180 247
rect 1200 227 1220 247
rect 1240 227 1260 247
rect 1280 227 1300 247
rect 1320 227 1340 247
rect 1360 227 1380 247
rect 1400 227 1420 247
rect 1440 227 1460 247
rect 1480 227 1500 247
rect 1520 227 1540 247
rect 1560 227 1580 247
rect 1600 227 1620 247
rect 1640 227 1660 247
rect 1680 227 1700 247
rect 1720 227 1740 247
rect 1760 227 1780 247
rect 1800 227 1820 247
rect 1840 227 1860 247
rect 1880 227 1900 247
rect 1920 227 1940 247
rect 1960 227 1980 247
rect 2000 227 2020 247
rect 2040 227 2060 247
rect 2080 227 2100 247
rect 2120 227 2140 247
rect 2160 227 2180 247
rect 2200 227 2220 247
rect 2240 227 2260 247
rect 2280 227 2300 247
rect 2320 227 2340 247
rect 2360 227 2380 247
rect 2400 227 2420 247
rect 2440 227 2460 247
rect 2480 227 2500 247
rect 2520 227 2540 247
rect 2560 227 2580 247
rect 2600 227 2620 247
rect 2640 227 2660 247
rect 200 145 220 165
rect 240 145 260 165
rect 280 145 300 165
rect 320 145 340 165
rect 360 145 380 165
rect 400 145 420 165
rect 440 145 460 165
rect 480 145 500 165
rect 520 145 540 165
rect 560 145 580 165
rect 600 145 620 165
rect 640 145 660 165
rect 680 145 700 165
rect 720 145 740 165
rect 760 145 780 165
rect 800 145 820 165
rect 840 145 860 165
rect 880 145 900 165
rect 920 145 940 165
rect 960 145 980 165
rect 1000 145 1020 165
rect 1040 145 1060 165
rect 1080 145 1100 165
rect 1120 145 1140 165
rect 1160 145 1180 165
rect 1200 145 1220 165
rect 1240 145 1260 165
rect 1280 145 1300 165
rect 1320 145 1340 165
rect 1360 145 1380 165
rect 1400 145 1420 165
rect 1440 145 1460 165
rect 1480 145 1500 165
rect 1520 145 1540 165
rect 1560 145 1580 165
rect 1600 145 1620 165
rect 1640 145 1660 165
rect 1680 145 1700 165
rect 1720 145 1740 165
rect 1760 145 1780 165
rect 1800 145 1820 165
rect 1840 145 1860 165
rect 1880 145 1900 165
rect 1920 145 1940 165
rect 1960 145 1980 165
rect 2000 145 2020 165
rect 2040 145 2060 165
rect 2080 145 2100 165
rect 2120 145 2140 165
rect 2160 145 2180 165
rect 2200 145 2220 165
rect 2240 145 2260 165
rect 2280 145 2300 165
rect 2320 145 2340 165
rect 2360 145 2380 165
rect 2400 145 2420 165
rect 2440 145 2460 165
rect 2480 145 2500 165
rect 2520 145 2540 165
rect 2560 145 2580 165
rect 2600 145 2620 165
rect 2640 145 2660 165
rect 120 -70 140 -50
rect 160 -70 180 -50
rect 200 -70 220 -50
rect 240 -70 260 -50
rect 280 -70 300 -50
rect 320 -70 340 -50
rect 360 -70 380 -50
rect 400 -70 420 -50
rect 440 -70 460 -50
rect 480 -70 500 -50
rect 520 -70 540 -50
rect 560 -70 580 -50
rect 600 -70 620 -50
rect 640 -70 660 -50
rect 680 -70 700 -50
rect 720 -70 740 -50
rect 760 -70 780 -50
rect 800 -70 820 -50
rect 840 -70 860 -50
rect 880 -70 900 -50
rect 920 -70 940 -50
rect 960 -70 980 -50
rect 1000 -70 1020 -50
rect 1040 -70 1060 -50
rect 1080 -70 1100 -50
rect 1120 -70 1140 -50
rect 1160 -70 1180 -50
rect 1200 -70 1220 -50
rect 1240 -70 1260 -50
rect 1280 -70 1300 -50
rect 1320 -70 1340 -50
rect 1360 -70 1380 -50
rect 1400 -70 1420 -50
rect 1440 -70 1460 -50
rect 1480 -70 1500 -50
rect 1520 -70 1540 -50
rect 1560 -70 1580 -50
rect 1600 -70 1620 -50
rect 1640 -70 1660 -50
rect 1680 -70 1700 -50
rect 1720 -70 1740 -50
rect 1760 -70 1780 -50
rect 1800 -70 1820 -50
rect 1840 -70 1860 -50
rect 1880 -70 1900 -50
rect 1920 -70 1940 -50
rect 1960 -70 1980 -50
rect 2000 -70 2020 -50
rect 2040 -70 2060 -50
rect 2080 -70 2100 -50
rect 2120 -70 2140 -50
rect 2160 -70 2180 -50
rect 2200 -70 2220 -50
rect 2240 -70 2260 -50
rect 2280 -70 2300 -50
rect 2320 -70 2340 -50
rect 2360 -70 2380 -50
rect 2400 -70 2420 -50
rect 2440 -70 2460 -50
rect 2480 -70 2500 -50
rect 2520 -70 2540 -50
rect 2560 -70 2590 -50
rect 120 -165 140 -145
rect 160 -165 180 -145
rect 200 -165 220 -145
rect 240 -165 260 -145
rect 280 -165 300 -145
rect 320 -165 340 -145
rect 360 -165 380 -145
rect 400 -165 420 -145
rect 440 -165 460 -145
rect 480 -165 500 -145
rect 520 -165 540 -145
rect 560 -165 580 -145
rect 600 -165 620 -145
rect 640 -165 660 -145
rect 680 -165 700 -145
rect 720 -165 740 -145
rect 760 -165 780 -145
rect 800 -165 820 -145
rect 840 -165 860 -145
rect 880 -165 900 -145
rect 920 -165 940 -145
rect 960 -165 980 -145
rect 1000 -165 1020 -145
rect 1040 -165 1060 -145
rect 1080 -165 1100 -145
rect 1120 -165 1140 -145
rect 1160 -165 1180 -145
rect 1200 -165 1220 -145
rect 1240 -165 1260 -145
rect 1280 -165 1300 -145
rect 1320 -165 1340 -145
rect 1360 -165 1380 -145
rect 1400 -165 1420 -145
rect 1440 -165 1460 -145
rect 1480 -165 1500 -145
rect 1520 -165 1540 -145
rect 1560 -165 1580 -145
rect 1600 -165 1620 -145
rect 1640 -165 1660 -145
rect 1680 -165 1700 -145
rect 1720 -165 1740 -145
rect 1760 -165 1780 -145
rect 1800 -165 1820 -145
rect 1840 -165 1860 -145
rect 1880 -165 1900 -145
rect 1920 -165 1940 -145
rect 1960 -165 1980 -145
rect 2000 -165 2020 -145
rect 2040 -165 2060 -145
rect 2080 -165 2100 -145
rect 2120 -165 2140 -145
rect 2160 -165 2180 -145
rect 2200 -165 2220 -145
rect 2240 -165 2260 -145
rect 2280 -165 2300 -145
rect 2320 -165 2340 -145
rect 2360 -165 2380 -145
rect 2400 -165 2420 -145
rect 2440 -165 2460 -145
rect 2480 -165 2500 -145
rect 2520 -165 2540 -145
rect 2560 -165 2590 -145
rect 120 -260 140 -240
rect 160 -260 180 -240
rect 200 -260 220 -240
rect 240 -260 260 -240
rect 280 -260 300 -240
rect 320 -260 340 -240
rect 360 -260 380 -240
rect 400 -260 420 -240
rect 440 -260 460 -240
rect 480 -260 500 -240
rect 520 -260 540 -240
rect 560 -260 580 -240
rect 600 -260 620 -240
rect 640 -260 660 -240
rect 680 -260 700 -240
rect 720 -260 740 -240
rect 760 -260 780 -240
rect 800 -260 820 -240
rect 840 -260 860 -240
rect 880 -260 900 -240
rect 920 -260 940 -240
rect 960 -260 980 -240
rect 1000 -260 1020 -240
rect 1040 -260 1060 -240
rect 1080 -260 1100 -240
rect 1120 -260 1140 -240
rect 1160 -260 1180 -240
rect 1200 -260 1220 -240
rect 1240 -260 1260 -240
rect 1280 -260 1300 -240
rect 1320 -260 1340 -240
rect 1360 -260 1380 -240
rect 1400 -260 1420 -240
rect 1440 -260 1460 -240
rect 1480 -260 1500 -240
rect 1520 -260 1540 -240
rect 1560 -260 1580 -240
rect 1600 -260 1620 -240
rect 1640 -260 1660 -240
rect 1680 -260 1700 -240
rect 1720 -260 1740 -240
rect 1760 -260 1780 -240
rect 1800 -260 1820 -240
rect 1840 -260 1860 -240
rect 1880 -260 1900 -240
rect 1920 -260 1940 -240
rect 1960 -260 1980 -240
rect 2000 -260 2020 -240
rect 2040 -260 2060 -240
rect 2080 -260 2100 -240
rect 2120 -260 2140 -240
rect 2160 -260 2180 -240
rect 2200 -260 2220 -240
rect 2240 -260 2260 -240
rect 2280 -260 2300 -240
rect 2320 -260 2340 -240
rect 2360 -260 2380 -240
rect 2400 -260 2420 -240
rect 2440 -260 2460 -240
rect 2480 -260 2500 -240
rect 2520 -260 2540 -240
rect 2560 -260 2590 -240
rect 120 -355 140 -335
rect 160 -355 180 -335
rect 200 -355 220 -335
rect 240 -355 260 -335
rect 280 -355 300 -335
rect 320 -355 340 -335
rect 360 -355 380 -335
rect 400 -355 420 -335
rect 440 -355 460 -335
rect 480 -355 500 -335
rect 520 -355 540 -335
rect 560 -355 580 -335
rect 600 -355 620 -335
rect 640 -355 660 -335
rect 680 -355 700 -335
rect 720 -355 740 -335
rect 760 -355 780 -335
rect 800 -355 820 -335
rect 840 -355 860 -335
rect 880 -355 900 -335
rect 920 -355 940 -335
rect 960 -355 980 -335
rect 1000 -355 1020 -335
rect 1040 -355 1060 -335
rect 1080 -355 1100 -335
rect 1120 -355 1140 -335
rect 1160 -355 1180 -335
rect 1200 -355 1220 -335
rect 1240 -355 1260 -335
rect 1280 -355 1300 -335
rect 1320 -355 1340 -335
rect 1360 -355 1380 -335
rect 1400 -355 1420 -335
rect 1440 -355 1460 -335
rect 1480 -355 1500 -335
rect 1520 -355 1540 -335
rect 1560 -355 1580 -335
rect 1600 -355 1620 -335
rect 1640 -355 1660 -335
rect 1680 -355 1700 -335
rect 1720 -355 1740 -335
rect 1760 -355 1780 -335
rect 1800 -355 1820 -335
rect 1840 -355 1860 -335
rect 1880 -355 1900 -335
rect 1920 -355 1940 -335
rect 1960 -355 1980 -335
rect 2000 -355 2020 -335
rect 2040 -355 2060 -335
rect 2080 -355 2100 -335
rect 2120 -355 2140 -335
rect 2160 -355 2180 -335
rect 2200 -355 2220 -335
rect 2240 -355 2260 -335
rect 2280 -355 2300 -335
rect 2320 -355 2340 -335
rect 2360 -355 2380 -335
rect 2400 -355 2420 -335
rect 2440 -355 2460 -335
rect 2480 -355 2500 -335
rect 2520 -355 2540 -335
rect 2560 -355 2590 -335
rect 120 -450 140 -430
rect 160 -450 180 -430
rect 200 -450 220 -430
rect 240 -450 260 -430
rect 280 -450 300 -430
rect 320 -450 340 -430
rect 360 -450 380 -430
rect 400 -450 420 -430
rect 440 -450 460 -430
rect 480 -450 500 -430
rect 520 -450 540 -430
rect 560 -450 580 -430
rect 600 -450 620 -430
rect 640 -450 660 -430
rect 680 -450 700 -430
rect 720 -450 740 -430
rect 760 -450 780 -430
rect 800 -450 820 -430
rect 840 -450 860 -430
rect 880 -450 900 -430
rect 920 -450 940 -430
rect 960 -450 980 -430
rect 1000 -450 1020 -430
rect 1040 -450 1060 -430
rect 1080 -450 1100 -430
rect 1120 -450 1140 -430
rect 1160 -450 1180 -430
rect 1200 -450 1220 -430
rect 1240 -450 1260 -430
rect 1280 -450 1300 -430
rect 1320 -450 1340 -430
rect 1360 -450 1380 -430
rect 1400 -450 1420 -430
rect 1440 -450 1460 -430
rect 1480 -450 1500 -430
rect 1520 -450 1540 -430
rect 1560 -450 1580 -430
rect 1600 -450 1620 -430
rect 1640 -450 1660 -430
rect 1680 -450 1700 -430
rect 1720 -450 1740 -430
rect 1760 -450 1780 -430
rect 1800 -450 1820 -430
rect 1840 -450 1860 -430
rect 1880 -450 1900 -430
rect 1920 -450 1940 -430
rect 1960 -450 1980 -430
rect 2000 -450 2020 -430
rect 2040 -450 2060 -430
rect 2080 -450 2100 -430
rect 2120 -450 2140 -430
rect 2160 -450 2180 -430
rect 2200 -450 2220 -430
rect 2240 -450 2260 -430
rect 2280 -450 2300 -430
rect 2320 -450 2340 -430
rect 2360 -450 2380 -430
rect 2400 -450 2420 -430
rect 2440 -450 2460 -430
rect 2480 -450 2500 -430
rect 2520 -450 2540 -430
rect 2560 -450 2590 -430
rect 120 -545 140 -525
rect 160 -545 180 -525
rect 200 -545 220 -525
rect 240 -545 260 -525
rect 280 -545 300 -525
rect 320 -545 340 -525
rect 360 -545 380 -525
rect 400 -545 420 -525
rect 440 -545 460 -525
rect 480 -545 500 -525
rect 520 -545 540 -525
rect 560 -545 580 -525
rect 600 -545 620 -525
rect 640 -545 660 -525
rect 680 -545 700 -525
rect 720 -545 740 -525
rect 760 -545 780 -525
rect 800 -545 820 -525
rect 840 -545 860 -525
rect 880 -545 900 -525
rect 920 -545 940 -525
rect 960 -545 980 -525
rect 1000 -545 1020 -525
rect 1040 -545 1060 -525
rect 1080 -545 1100 -525
rect 1120 -545 1140 -525
rect 1160 -545 1180 -525
rect 1200 -545 1220 -525
rect 1240 -545 1260 -525
rect 1280 -545 1300 -525
rect 1320 -545 1340 -525
rect 1360 -545 1380 -525
rect 1400 -545 1420 -525
rect 1440 -545 1460 -525
rect 1480 -545 1500 -525
rect 1520 -545 1540 -525
rect 1560 -545 1580 -525
rect 1600 -545 1620 -525
rect 1640 -545 1660 -525
rect 1680 -545 1700 -525
rect 1720 -545 1740 -525
rect 1760 -545 1780 -525
rect 1800 -545 1820 -525
rect 1840 -545 1860 -525
rect 1880 -545 1900 -525
rect 1920 -545 1940 -525
rect 1960 -545 1980 -525
rect 2000 -545 2020 -525
rect 2040 -545 2060 -525
rect 2080 -545 2100 -525
rect 2120 -545 2140 -525
rect 2160 -545 2180 -525
rect 2200 -545 2220 -525
rect 2240 -545 2260 -525
rect 2280 -545 2300 -525
rect 2320 -545 2340 -525
rect 2360 -545 2380 -525
rect 2400 -545 2420 -525
rect 2440 -545 2460 -525
rect 2480 -545 2500 -525
rect 2520 -545 2540 -525
rect 2560 -545 2590 -525
rect 120 -640 140 -620
rect 160 -640 180 -620
rect 200 -640 220 -620
rect 240 -640 260 -620
rect 280 -640 300 -620
rect 320 -640 340 -620
rect 360 -640 380 -620
rect 400 -640 420 -620
rect 440 -640 460 -620
rect 480 -640 500 -620
rect 520 -640 540 -620
rect 560 -640 580 -620
rect 600 -640 620 -620
rect 640 -640 660 -620
rect 680 -640 700 -620
rect 720 -640 740 -620
rect 760 -640 780 -620
rect 800 -640 820 -620
rect 840 -640 860 -620
rect 880 -640 900 -620
rect 920 -640 940 -620
rect 960 -640 980 -620
rect 1000 -640 1020 -620
rect 1040 -640 1060 -620
rect 1080 -640 1100 -620
rect 1120 -640 1140 -620
rect 1160 -640 1180 -620
rect 1200 -640 1220 -620
rect 1240 -640 1260 -620
rect 1280 -640 1300 -620
rect 1320 -640 1340 -620
rect 1360 -640 1380 -620
rect 1400 -640 1420 -620
rect 1440 -640 1460 -620
rect 1480 -640 1500 -620
rect 1520 -640 1540 -620
rect 1560 -640 1580 -620
rect 1600 -640 1620 -620
rect 1640 -640 1660 -620
rect 1680 -640 1700 -620
rect 1720 -640 1740 -620
rect 1760 -640 1780 -620
rect 1800 -640 1820 -620
rect 1840 -640 1860 -620
rect 1880 -640 1900 -620
rect 1920 -640 1940 -620
rect 1960 -640 1980 -620
rect 2000 -640 2020 -620
rect 2040 -640 2060 -620
rect 2080 -640 2100 -620
rect 2120 -640 2140 -620
rect 2160 -640 2180 -620
rect 2200 -640 2220 -620
rect 2240 -640 2260 -620
rect 2280 -640 2300 -620
rect 2320 -640 2340 -620
rect 2360 -640 2380 -620
rect 2400 -640 2420 -620
rect 2440 -640 2460 -620
rect 2480 -640 2500 -620
rect 2520 -640 2540 -620
rect 2560 -640 2590 -620
rect 120 -735 140 -715
rect 160 -735 180 -715
rect 200 -735 220 -715
rect 240 -735 260 -715
rect 280 -735 300 -715
rect 320 -735 340 -715
rect 360 -735 380 -715
rect 400 -735 420 -715
rect 440 -735 460 -715
rect 480 -735 500 -715
rect 520 -735 540 -715
rect 560 -735 580 -715
rect 600 -735 620 -715
rect 640 -735 660 -715
rect 680 -735 700 -715
rect 720 -735 740 -715
rect 760 -735 780 -715
rect 800 -735 820 -715
rect 840 -735 860 -715
rect 880 -735 900 -715
rect 920 -735 940 -715
rect 960 -735 980 -715
rect 1000 -735 1020 -715
rect 1040 -735 1060 -715
rect 1080 -735 1100 -715
rect 1120 -735 1140 -715
rect 1160 -735 1180 -715
rect 1200 -735 1220 -715
rect 1240 -735 1260 -715
rect 1280 -735 1300 -715
rect 1320 -735 1340 -715
rect 1360 -735 1380 -715
rect 1400 -735 1420 -715
rect 1440 -735 1460 -715
rect 1480 -735 1500 -715
rect 1520 -735 1540 -715
rect 1560 -735 1580 -715
rect 1600 -735 1620 -715
rect 1640 -735 1660 -715
rect 1680 -735 1700 -715
rect 1720 -735 1740 -715
rect 1760 -735 1780 -715
rect 1800 -735 1820 -715
rect 1840 -735 1860 -715
rect 1880 -735 1900 -715
rect 1920 -735 1940 -715
rect 1960 -735 1980 -715
rect 2000 -735 2020 -715
rect 2040 -735 2060 -715
rect 2080 -735 2100 -715
rect 2120 -735 2140 -715
rect 2160 -735 2180 -715
rect 2200 -735 2220 -715
rect 2240 -735 2260 -715
rect 2280 -735 2300 -715
rect 2320 -735 2340 -715
rect 2360 -735 2380 -715
rect 2400 -735 2420 -715
rect 2440 -735 2460 -715
rect 2480 -735 2500 -715
rect 2520 -735 2540 -715
rect 2560 -735 2590 -715
rect 120 -830 140 -810
rect 160 -830 180 -810
rect 200 -830 220 -810
rect 240 -830 260 -810
rect 280 -830 300 -810
rect 320 -830 340 -810
rect 360 -830 380 -810
rect 400 -830 420 -810
rect 440 -830 460 -810
rect 480 -830 500 -810
rect 520 -830 540 -810
rect 560 -830 580 -810
rect 600 -830 620 -810
rect 640 -830 660 -810
rect 680 -830 700 -810
rect 720 -830 740 -810
rect 760 -830 780 -810
rect 800 -830 820 -810
rect 840 -830 860 -810
rect 880 -830 900 -810
rect 920 -830 940 -810
rect 960 -830 980 -810
rect 1000 -830 1020 -810
rect 1040 -830 1060 -810
rect 1080 -830 1100 -810
rect 1120 -830 1140 -810
rect 1160 -830 1180 -810
rect 1200 -830 1220 -810
rect 1240 -830 1260 -810
rect 1280 -830 1300 -810
rect 1320 -830 1340 -810
rect 1360 -830 1380 -810
rect 1400 -830 1420 -810
rect 1440 -830 1460 -810
rect 1480 -830 1500 -810
rect 1520 -830 1540 -810
rect 1560 -830 1580 -810
rect 1600 -830 1620 -810
rect 1640 -830 1660 -810
rect 1680 -830 1700 -810
rect 1720 -830 1740 -810
rect 1760 -830 1780 -810
rect 1800 -830 1820 -810
rect 1840 -830 1860 -810
rect 1880 -830 1900 -810
rect 1920 -830 1940 -810
rect 1960 -830 1980 -810
rect 2000 -830 2020 -810
rect 2040 -830 2060 -810
rect 2080 -830 2100 -810
rect 2120 -830 2140 -810
rect 2160 -830 2180 -810
rect 2200 -830 2220 -810
rect 2240 -830 2260 -810
rect 2280 -830 2300 -810
rect 2320 -830 2340 -810
rect 2360 -830 2380 -810
rect 2400 -830 2420 -810
rect 2440 -830 2460 -810
rect 2480 -830 2500 -810
rect 2520 -830 2540 -810
rect 2560 -830 2590 -810
rect 120 -925 140 -905
rect 160 -925 180 -905
rect 200 -925 220 -905
rect 240 -925 260 -905
rect 280 -925 300 -905
rect 320 -925 340 -905
rect 360 -925 380 -905
rect 400 -925 420 -905
rect 440 -925 460 -905
rect 480 -925 500 -905
rect 520 -925 540 -905
rect 560 -925 580 -905
rect 600 -925 620 -905
rect 640 -925 660 -905
rect 680 -925 700 -905
rect 720 -925 740 -905
rect 760 -925 780 -905
rect 800 -925 820 -905
rect 840 -925 860 -905
rect 880 -925 900 -905
rect 920 -925 940 -905
rect 960 -925 980 -905
rect 1000 -925 1020 -905
rect 1040 -925 1060 -905
rect 1080 -925 1100 -905
rect 1120 -925 1140 -905
rect 1160 -925 1180 -905
rect 1200 -925 1220 -905
rect 1240 -925 1260 -905
rect 1280 -925 1300 -905
rect 1320 -925 1340 -905
rect 1360 -925 1380 -905
rect 1400 -925 1420 -905
rect 1440 -925 1460 -905
rect 1480 -925 1500 -905
rect 1520 -925 1540 -905
rect 1560 -925 1580 -905
rect 1600 -925 1620 -905
rect 1640 -925 1660 -905
rect 1680 -925 1700 -905
rect 1720 -925 1740 -905
rect 1760 -925 1780 -905
rect 1800 -925 1820 -905
rect 1840 -925 1860 -905
rect 1880 -925 1900 -905
rect 1920 -925 1940 -905
rect 1960 -925 1980 -905
rect 2000 -925 2020 -905
rect 2040 -925 2060 -905
rect 2080 -925 2100 -905
rect 2120 -925 2140 -905
rect 2160 -925 2180 -905
rect 2200 -925 2220 -905
rect 2240 -925 2260 -905
rect 2280 -925 2300 -905
rect 2320 -925 2340 -905
rect 2360 -925 2380 -905
rect 2400 -925 2420 -905
rect 2440 -925 2460 -905
rect 2480 -925 2500 -905
rect 2520 -925 2540 -905
rect 2560 -925 2590 -905
rect 120 -1020 140 -1000
rect 160 -1020 180 -1000
rect 200 -1020 220 -1000
rect 240 -1020 260 -1000
rect 280 -1020 300 -1000
rect 320 -1020 340 -1000
rect 360 -1020 380 -1000
rect 400 -1020 420 -1000
rect 440 -1020 460 -1000
rect 480 -1020 500 -1000
rect 520 -1020 540 -1000
rect 560 -1020 580 -1000
rect 600 -1020 620 -1000
rect 640 -1020 660 -1000
rect 680 -1020 700 -1000
rect 720 -1020 740 -1000
rect 760 -1020 780 -1000
rect 800 -1020 820 -1000
rect 840 -1020 860 -1000
rect 880 -1020 900 -1000
rect 920 -1020 940 -1000
rect 960 -1020 980 -1000
rect 1000 -1020 1020 -1000
rect 1040 -1020 1060 -1000
rect 1080 -1020 1100 -1000
rect 1120 -1020 1140 -1000
rect 1160 -1020 1180 -1000
rect 1200 -1020 1220 -1000
rect 1240 -1020 1260 -1000
rect 1280 -1020 1300 -1000
rect 1320 -1020 1340 -1000
rect 1360 -1020 1380 -1000
rect 1400 -1020 1420 -1000
rect 1440 -1020 1460 -1000
rect 1480 -1020 1500 -1000
rect 1520 -1020 1540 -1000
rect 1560 -1020 1580 -1000
rect 1600 -1020 1620 -1000
rect 1640 -1020 1660 -1000
rect 1680 -1020 1700 -1000
rect 1720 -1020 1740 -1000
rect 1760 -1020 1780 -1000
rect 1800 -1020 1820 -1000
rect 1840 -1020 1860 -1000
rect 1880 -1020 1900 -1000
rect 1920 -1020 1940 -1000
rect 1960 -1020 1980 -1000
rect 2000 -1020 2020 -1000
rect 2040 -1020 2060 -1000
rect 2080 -1020 2100 -1000
rect 2120 -1020 2140 -1000
rect 2160 -1020 2180 -1000
rect 2200 -1020 2220 -1000
rect 2240 -1020 2260 -1000
rect 2280 -1020 2300 -1000
rect 2320 -1020 2340 -1000
rect 2360 -1020 2380 -1000
rect 2400 -1020 2420 -1000
rect 2440 -1020 2460 -1000
rect 2480 -1020 2500 -1000
rect 2520 -1020 2540 -1000
rect 2560 -1020 2590 -1000
rect 120 -1115 140 -1095
rect 160 -1115 180 -1095
rect 200 -1115 220 -1095
rect 240 -1115 260 -1095
rect 280 -1115 300 -1095
rect 320 -1115 340 -1095
rect 360 -1115 380 -1095
rect 400 -1115 420 -1095
rect 440 -1115 460 -1095
rect 480 -1115 500 -1095
rect 520 -1115 540 -1095
rect 560 -1115 580 -1095
rect 600 -1115 620 -1095
rect 640 -1115 660 -1095
rect 680 -1115 700 -1095
rect 720 -1115 740 -1095
rect 760 -1115 780 -1095
rect 800 -1115 820 -1095
rect 840 -1115 860 -1095
rect 880 -1115 900 -1095
rect 920 -1115 940 -1095
rect 960 -1115 980 -1095
rect 1000 -1115 1020 -1095
rect 1040 -1115 1060 -1095
rect 1080 -1115 1100 -1095
rect 1120 -1115 1140 -1095
rect 1160 -1115 1180 -1095
rect 1200 -1115 1220 -1095
rect 1240 -1115 1260 -1095
rect 1280 -1115 1300 -1095
rect 1320 -1115 1340 -1095
rect 1360 -1115 1380 -1095
rect 1400 -1115 1420 -1095
rect 1440 -1115 1460 -1095
rect 1480 -1115 1500 -1095
rect 1520 -1115 1540 -1095
rect 1560 -1115 1580 -1095
rect 1600 -1115 1620 -1095
rect 1640 -1115 1660 -1095
rect 1680 -1115 1700 -1095
rect 1720 -1115 1740 -1095
rect 1760 -1115 1780 -1095
rect 1800 -1115 1820 -1095
rect 1840 -1115 1860 -1095
rect 1880 -1115 1900 -1095
rect 1920 -1115 1940 -1095
rect 1960 -1115 1980 -1095
rect 2000 -1115 2020 -1095
rect 2040 -1115 2060 -1095
rect 2080 -1115 2100 -1095
rect 2120 -1115 2140 -1095
rect 2160 -1115 2180 -1095
rect 2200 -1115 2220 -1095
rect 2240 -1115 2260 -1095
rect 2280 -1115 2300 -1095
rect 2320 -1115 2340 -1095
rect 2360 -1115 2380 -1095
rect 2400 -1115 2420 -1095
rect 2440 -1115 2460 -1095
rect 2480 -1115 2500 -1095
rect 2520 -1115 2540 -1095
rect 2560 -1115 2590 -1095
rect 120 -1210 140 -1190
rect 160 -1210 180 -1190
rect 200 -1210 220 -1190
rect 240 -1210 260 -1190
rect 280 -1210 300 -1190
rect 320 -1210 340 -1190
rect 360 -1210 380 -1190
rect 400 -1210 420 -1190
rect 440 -1210 460 -1190
rect 480 -1210 500 -1190
rect 520 -1210 540 -1190
rect 560 -1210 580 -1190
rect 600 -1210 620 -1190
rect 640 -1210 660 -1190
rect 680 -1210 700 -1190
rect 720 -1210 740 -1190
rect 760 -1210 780 -1190
rect 800 -1210 820 -1190
rect 840 -1210 860 -1190
rect 880 -1210 900 -1190
rect 920 -1210 940 -1190
rect 960 -1210 980 -1190
rect 1000 -1210 1020 -1190
rect 1040 -1210 1060 -1190
rect 1080 -1210 1100 -1190
rect 1120 -1210 1140 -1190
rect 1160 -1210 1180 -1190
rect 1200 -1210 1220 -1190
rect 1240 -1210 1260 -1190
rect 1280 -1210 1300 -1190
rect 1320 -1210 1340 -1190
rect 1360 -1210 1380 -1190
rect 1400 -1210 1420 -1190
rect 1440 -1210 1460 -1190
rect 1480 -1210 1500 -1190
rect 1520 -1210 1540 -1190
rect 1560 -1210 1580 -1190
rect 1600 -1210 1620 -1190
rect 1640 -1210 1660 -1190
rect 1680 -1210 1700 -1190
rect 1720 -1210 1740 -1190
rect 1760 -1210 1780 -1190
rect 1800 -1210 1820 -1190
rect 1840 -1210 1860 -1190
rect 1880 -1210 1900 -1190
rect 1920 -1210 1940 -1190
rect 1960 -1210 1980 -1190
rect 2000 -1210 2020 -1190
rect 2040 -1210 2060 -1190
rect 2080 -1210 2100 -1190
rect 2120 -1210 2140 -1190
rect 2160 -1210 2180 -1190
rect 2200 -1210 2220 -1190
rect 2240 -1210 2260 -1190
rect 2280 -1210 2300 -1190
rect 2320 -1210 2340 -1190
rect 2360 -1210 2380 -1190
rect 2400 -1210 2420 -1190
rect 2440 -1210 2460 -1190
rect 2480 -1210 2500 -1190
rect 2520 -1210 2540 -1190
rect 2560 -1210 2590 -1190
rect 120 -1305 140 -1285
rect 160 -1305 180 -1285
rect 200 -1305 220 -1285
rect 240 -1305 260 -1285
rect 280 -1305 300 -1285
rect 320 -1305 340 -1285
rect 360 -1305 380 -1285
rect 400 -1305 420 -1285
rect 440 -1305 460 -1285
rect 480 -1305 500 -1285
rect 520 -1305 540 -1285
rect 560 -1305 580 -1285
rect 600 -1305 620 -1285
rect 640 -1305 660 -1285
rect 680 -1305 700 -1285
rect 720 -1305 740 -1285
rect 760 -1305 780 -1285
rect 800 -1305 820 -1285
rect 840 -1305 860 -1285
rect 880 -1305 900 -1285
rect 920 -1305 940 -1285
rect 960 -1305 980 -1285
rect 1000 -1305 1020 -1285
rect 1040 -1305 1060 -1285
rect 1080 -1305 1100 -1285
rect 1120 -1305 1140 -1285
rect 1160 -1305 1180 -1285
rect 1200 -1305 1220 -1285
rect 1240 -1305 1260 -1285
rect 1280 -1305 1300 -1285
rect 1320 -1305 1340 -1285
rect 1360 -1305 1380 -1285
rect 1400 -1305 1420 -1285
rect 1440 -1305 1460 -1285
rect 1480 -1305 1500 -1285
rect 1520 -1305 1540 -1285
rect 1560 -1305 1580 -1285
rect 1600 -1305 1620 -1285
rect 1640 -1305 1660 -1285
rect 1680 -1305 1700 -1285
rect 1720 -1305 1740 -1285
rect 1760 -1305 1780 -1285
rect 1800 -1305 1820 -1285
rect 1840 -1305 1860 -1285
rect 1880 -1305 1900 -1285
rect 1920 -1305 1940 -1285
rect 1960 -1305 1980 -1285
rect 2000 -1305 2020 -1285
rect 2040 -1305 2060 -1285
rect 2080 -1305 2100 -1285
rect 2120 -1305 2140 -1285
rect 2160 -1305 2180 -1285
rect 2200 -1305 2220 -1285
rect 2240 -1305 2260 -1285
rect 2280 -1305 2300 -1285
rect 2320 -1305 2340 -1285
rect 2360 -1305 2380 -1285
rect 2400 -1305 2420 -1285
rect 2440 -1305 2460 -1285
rect 2480 -1305 2500 -1285
rect 2520 -1305 2540 -1285
rect 2560 -1305 2590 -1285
rect 120 -1400 140 -1380
rect 160 -1400 180 -1380
rect 200 -1400 220 -1380
rect 240 -1400 260 -1380
rect 280 -1400 300 -1380
rect 320 -1400 340 -1380
rect 360 -1400 380 -1380
rect 400 -1400 420 -1380
rect 440 -1400 460 -1380
rect 480 -1400 500 -1380
rect 520 -1400 540 -1380
rect 560 -1400 580 -1380
rect 600 -1400 620 -1380
rect 640 -1400 660 -1380
rect 680 -1400 700 -1380
rect 720 -1400 740 -1380
rect 760 -1400 780 -1380
rect 800 -1400 820 -1380
rect 840 -1400 860 -1380
rect 880 -1400 900 -1380
rect 920 -1400 940 -1380
rect 960 -1400 980 -1380
rect 1000 -1400 1020 -1380
rect 1040 -1400 1060 -1380
rect 1080 -1400 1100 -1380
rect 1120 -1400 1140 -1380
rect 1160 -1400 1180 -1380
rect 1200 -1400 1220 -1380
rect 1240 -1400 1260 -1380
rect 1280 -1400 1300 -1380
rect 1320 -1400 1340 -1380
rect 1360 -1400 1380 -1380
rect 1400 -1400 1420 -1380
rect 1440 -1400 1460 -1380
rect 1480 -1400 1500 -1380
rect 1520 -1400 1540 -1380
rect 1560 -1400 1580 -1380
rect 1600 -1400 1620 -1380
rect 1640 -1400 1660 -1380
rect 1680 -1400 1700 -1380
rect 1720 -1400 1740 -1380
rect 1760 -1400 1780 -1380
rect 1800 -1400 1820 -1380
rect 1840 -1400 1860 -1380
rect 1880 -1400 1900 -1380
rect 1920 -1400 1940 -1380
rect 1960 -1400 1980 -1380
rect 2000 -1400 2020 -1380
rect 2040 -1400 2060 -1380
rect 2080 -1400 2100 -1380
rect 2120 -1400 2140 -1380
rect 2160 -1400 2180 -1380
rect 2200 -1400 2220 -1380
rect 2240 -1400 2260 -1380
rect 2280 -1400 2300 -1380
rect 2320 -1400 2340 -1380
rect 2360 -1400 2380 -1380
rect 2400 -1400 2420 -1380
rect 2440 -1400 2460 -1380
rect 2480 -1400 2500 -1380
rect 2520 -1400 2540 -1380
rect 2560 -1400 2590 -1380
rect 120 -1495 140 -1475
rect 160 -1495 180 -1475
rect 200 -1495 220 -1475
rect 240 -1495 260 -1475
rect 280 -1495 300 -1475
rect 320 -1495 340 -1475
rect 360 -1495 380 -1475
rect 400 -1495 420 -1475
rect 440 -1495 460 -1475
rect 480 -1495 500 -1475
rect 520 -1495 540 -1475
rect 560 -1495 580 -1475
rect 600 -1495 620 -1475
rect 640 -1495 660 -1475
rect 680 -1495 700 -1475
rect 720 -1495 740 -1475
rect 760 -1495 780 -1475
rect 800 -1495 820 -1475
rect 840 -1495 860 -1475
rect 880 -1495 900 -1475
rect 920 -1495 940 -1475
rect 960 -1495 980 -1475
rect 1000 -1495 1020 -1475
rect 1040 -1495 1060 -1475
rect 1080 -1495 1100 -1475
rect 1120 -1495 1140 -1475
rect 1160 -1495 1180 -1475
rect 1200 -1495 1220 -1475
rect 1240 -1495 1260 -1475
rect 1280 -1495 1300 -1475
rect 1320 -1495 1340 -1475
rect 1360 -1495 1380 -1475
rect 1400 -1495 1420 -1475
rect 1440 -1495 1460 -1475
rect 1480 -1495 1500 -1475
rect 1520 -1495 1540 -1475
rect 1560 -1495 1580 -1475
rect 1600 -1495 1620 -1475
rect 1640 -1495 1660 -1475
rect 1680 -1495 1700 -1475
rect 1720 -1495 1740 -1475
rect 1760 -1495 1780 -1475
rect 1800 -1495 1820 -1475
rect 1840 -1495 1860 -1475
rect 1880 -1495 1900 -1475
rect 1920 -1495 1940 -1475
rect 1960 -1495 1980 -1475
rect 2000 -1495 2020 -1475
rect 2040 -1495 2060 -1475
rect 2080 -1495 2100 -1475
rect 2120 -1495 2140 -1475
rect 2160 -1495 2180 -1475
rect 2200 -1495 2220 -1475
rect 2240 -1495 2260 -1475
rect 2280 -1495 2300 -1475
rect 2320 -1495 2340 -1475
rect 2360 -1495 2380 -1475
rect 2400 -1495 2420 -1475
rect 2440 -1495 2460 -1475
rect 2480 -1495 2500 -1475
rect 2520 -1495 2540 -1475
rect 2560 -1495 2590 -1475
rect 120 -1590 140 -1570
rect 160 -1590 180 -1570
rect 200 -1590 220 -1570
rect 240 -1590 260 -1570
rect 280 -1590 300 -1570
rect 320 -1590 340 -1570
rect 360 -1590 380 -1570
rect 400 -1590 420 -1570
rect 440 -1590 460 -1570
rect 480 -1590 500 -1570
rect 520 -1590 540 -1570
rect 560 -1590 580 -1570
rect 600 -1590 620 -1570
rect 640 -1590 660 -1570
rect 680 -1590 700 -1570
rect 720 -1590 740 -1570
rect 760 -1590 780 -1570
rect 800 -1590 820 -1570
rect 840 -1590 860 -1570
rect 880 -1590 900 -1570
rect 920 -1590 940 -1570
rect 960 -1590 980 -1570
rect 1000 -1590 1020 -1570
rect 1040 -1590 1060 -1570
rect 1080 -1590 1100 -1570
rect 1120 -1590 1140 -1570
rect 1160 -1590 1180 -1570
rect 1200 -1590 1220 -1570
rect 1240 -1590 1260 -1570
rect 1280 -1590 1300 -1570
rect 1320 -1590 1340 -1570
rect 1360 -1590 1380 -1570
rect 1400 -1590 1420 -1570
rect 1440 -1590 1460 -1570
rect 1480 -1590 1500 -1570
rect 1520 -1590 1540 -1570
rect 1560 -1590 1580 -1570
rect 1600 -1590 1620 -1570
rect 1640 -1590 1660 -1570
rect 1680 -1590 1700 -1570
rect 1720 -1590 1740 -1570
rect 1760 -1590 1780 -1570
rect 1800 -1590 1820 -1570
rect 1840 -1590 1860 -1570
rect 1880 -1590 1900 -1570
rect 1920 -1590 1940 -1570
rect 1960 -1590 1980 -1570
rect 2000 -1590 2020 -1570
rect 2040 -1590 2060 -1570
rect 2080 -1590 2100 -1570
rect 2120 -1590 2140 -1570
rect 2160 -1590 2180 -1570
rect 2200 -1590 2220 -1570
rect 2240 -1590 2260 -1570
rect 2280 -1590 2300 -1570
rect 2320 -1590 2340 -1570
rect 2360 -1590 2380 -1570
rect 2400 -1590 2420 -1570
rect 2440 -1590 2460 -1570
rect 2480 -1590 2500 -1570
rect 2520 -1590 2540 -1570
rect 2560 -1590 2590 -1570
rect 120 -1685 140 -1665
rect 160 -1685 180 -1665
rect 200 -1685 220 -1665
rect 240 -1685 260 -1665
rect 280 -1685 300 -1665
rect 320 -1685 340 -1665
rect 360 -1685 380 -1665
rect 400 -1685 420 -1665
rect 440 -1685 460 -1665
rect 480 -1685 500 -1665
rect 520 -1685 540 -1665
rect 560 -1685 580 -1665
rect 600 -1685 620 -1665
rect 640 -1685 660 -1665
rect 680 -1685 700 -1665
rect 720 -1685 740 -1665
rect 760 -1685 780 -1665
rect 800 -1685 820 -1665
rect 840 -1685 860 -1665
rect 880 -1685 900 -1665
rect 920 -1685 940 -1665
rect 960 -1685 980 -1665
rect 1000 -1685 1020 -1665
rect 1040 -1685 1060 -1665
rect 1080 -1685 1100 -1665
rect 1120 -1685 1140 -1665
rect 1160 -1685 1180 -1665
rect 1200 -1685 1220 -1665
rect 1240 -1685 1260 -1665
rect 1280 -1685 1300 -1665
rect 1320 -1685 1340 -1665
rect 1360 -1685 1380 -1665
rect 1400 -1685 1420 -1665
rect 1440 -1685 1460 -1665
rect 1480 -1685 1500 -1665
rect 1520 -1685 1540 -1665
rect 1560 -1685 1580 -1665
rect 1600 -1685 1620 -1665
rect 1640 -1685 1660 -1665
rect 1680 -1685 1700 -1665
rect 1720 -1685 1740 -1665
rect 1760 -1685 1780 -1665
rect 1800 -1685 1820 -1665
rect 1840 -1685 1860 -1665
rect 1880 -1685 1900 -1665
rect 1920 -1685 1940 -1665
rect 1960 -1685 1980 -1665
rect 2000 -1685 2020 -1665
rect 2040 -1685 2060 -1665
rect 2080 -1685 2100 -1665
rect 2120 -1685 2140 -1665
rect 2160 -1685 2180 -1665
rect 2200 -1685 2220 -1665
rect 2240 -1685 2260 -1665
rect 2280 -1685 2300 -1665
rect 2320 -1685 2340 -1665
rect 2360 -1685 2380 -1665
rect 2400 -1685 2420 -1665
rect 2440 -1685 2460 -1665
rect 2480 -1685 2500 -1665
rect 2520 -1685 2540 -1665
rect 2560 -1685 2590 -1665
rect 120 -1780 140 -1760
rect 160 -1780 180 -1760
rect 200 -1780 220 -1760
rect 240 -1780 260 -1760
rect 280 -1780 300 -1760
rect 320 -1780 340 -1760
rect 360 -1780 380 -1760
rect 400 -1780 420 -1760
rect 440 -1780 460 -1760
rect 480 -1780 500 -1760
rect 520 -1780 540 -1760
rect 560 -1780 580 -1760
rect 600 -1780 620 -1760
rect 640 -1780 660 -1760
rect 680 -1780 700 -1760
rect 720 -1780 740 -1760
rect 760 -1780 780 -1760
rect 800 -1780 820 -1760
rect 840 -1780 860 -1760
rect 880 -1780 900 -1760
rect 920 -1780 940 -1760
rect 960 -1780 980 -1760
rect 1000 -1780 1020 -1760
rect 1040 -1780 1060 -1760
rect 1080 -1780 1100 -1760
rect 1120 -1780 1140 -1760
rect 1160 -1780 1180 -1760
rect 1200 -1780 1220 -1760
rect 1240 -1780 1260 -1760
rect 1280 -1780 1300 -1760
rect 1320 -1780 1340 -1760
rect 1360 -1780 1380 -1760
rect 1400 -1780 1420 -1760
rect 1440 -1780 1460 -1760
rect 1480 -1780 1500 -1760
rect 1520 -1780 1540 -1760
rect 1560 -1780 1580 -1760
rect 1600 -1780 1620 -1760
rect 1640 -1780 1660 -1760
rect 1680 -1780 1700 -1760
rect 1720 -1780 1740 -1760
rect 1760 -1780 1780 -1760
rect 1800 -1780 1820 -1760
rect 1840 -1780 1860 -1760
rect 1880 -1780 1900 -1760
rect 1920 -1780 1940 -1760
rect 1960 -1780 1980 -1760
rect 2000 -1780 2020 -1760
rect 2040 -1780 2060 -1760
rect 2080 -1780 2100 -1760
rect 2120 -1780 2140 -1760
rect 2160 -1780 2180 -1760
rect 2200 -1780 2220 -1760
rect 2240 -1780 2260 -1760
rect 2280 -1780 2300 -1760
rect 2320 -1780 2340 -1760
rect 2360 -1780 2380 -1760
rect 2400 -1780 2420 -1760
rect 2440 -1780 2460 -1760
rect 2480 -1780 2500 -1760
rect 2520 -1780 2540 -1760
rect 2560 -1780 2590 -1760
rect 120 -1875 140 -1855
rect 160 -1875 180 -1855
rect 200 -1875 220 -1855
rect 240 -1875 260 -1855
rect 280 -1875 300 -1855
rect 320 -1875 340 -1855
rect 360 -1875 380 -1855
rect 400 -1875 420 -1855
rect 440 -1875 460 -1855
rect 480 -1875 500 -1855
rect 520 -1875 540 -1855
rect 560 -1875 580 -1855
rect 600 -1875 620 -1855
rect 640 -1875 660 -1855
rect 680 -1875 700 -1855
rect 720 -1875 740 -1855
rect 760 -1875 780 -1855
rect 800 -1875 820 -1855
rect 840 -1875 860 -1855
rect 880 -1875 900 -1855
rect 920 -1875 940 -1855
rect 960 -1875 980 -1855
rect 1000 -1875 1020 -1855
rect 1040 -1875 1060 -1855
rect 1080 -1875 1100 -1855
rect 1120 -1875 1140 -1855
rect 1160 -1875 1180 -1855
rect 1200 -1875 1220 -1855
rect 1240 -1875 1260 -1855
rect 1280 -1875 1300 -1855
rect 1320 -1875 1340 -1855
rect 1360 -1875 1380 -1855
rect 1400 -1875 1420 -1855
rect 1440 -1875 1460 -1855
rect 1480 -1875 1500 -1855
rect 1520 -1875 1540 -1855
rect 1560 -1875 1580 -1855
rect 1600 -1875 1620 -1855
rect 1640 -1875 1660 -1855
rect 1680 -1875 1700 -1855
rect 1720 -1875 1740 -1855
rect 1760 -1875 1780 -1855
rect 1800 -1875 1820 -1855
rect 1840 -1875 1860 -1855
rect 1880 -1875 1900 -1855
rect 1920 -1875 1940 -1855
rect 1960 -1875 1980 -1855
rect 2000 -1875 2020 -1855
rect 2040 -1875 2060 -1855
rect 2080 -1875 2100 -1855
rect 2120 -1875 2140 -1855
rect 2160 -1875 2180 -1855
rect 2200 -1875 2220 -1855
rect 2240 -1875 2260 -1855
rect 2280 -1875 2300 -1855
rect 2320 -1875 2340 -1855
rect 2360 -1875 2380 -1855
rect 2400 -1875 2420 -1855
rect 2440 -1875 2460 -1855
rect 2480 -1875 2500 -1855
rect 2520 -1875 2540 -1855
rect 2560 -1875 2590 -1855
rect 120 -1970 140 -1950
rect 160 -1970 180 -1950
rect 200 -1970 220 -1950
rect 240 -1970 260 -1950
rect 280 -1970 300 -1950
rect 320 -1970 340 -1950
rect 360 -1970 380 -1950
rect 400 -1970 420 -1950
rect 440 -1970 460 -1950
rect 480 -1970 500 -1950
rect 520 -1970 540 -1950
rect 560 -1970 580 -1950
rect 600 -1970 620 -1950
rect 640 -1970 660 -1950
rect 680 -1970 700 -1950
rect 720 -1970 740 -1950
rect 760 -1970 780 -1950
rect 800 -1970 820 -1950
rect 840 -1970 860 -1950
rect 880 -1970 900 -1950
rect 920 -1970 940 -1950
rect 960 -1970 980 -1950
rect 1000 -1970 1020 -1950
rect 1040 -1970 1060 -1950
rect 1080 -1970 1100 -1950
rect 1120 -1970 1140 -1950
rect 1160 -1970 1180 -1950
rect 1200 -1970 1220 -1950
rect 1240 -1970 1260 -1950
rect 1280 -1970 1300 -1950
rect 1320 -1970 1340 -1950
rect 1360 -1970 1380 -1950
rect 1400 -1970 1420 -1950
rect 1440 -1970 1460 -1950
rect 1480 -1970 1500 -1950
rect 1520 -1970 1540 -1950
rect 1560 -1970 1580 -1950
rect 1600 -1970 1620 -1950
rect 1640 -1970 1660 -1950
rect 1680 -1970 1700 -1950
rect 1720 -1970 1740 -1950
rect 1760 -1970 1780 -1950
rect 1800 -1970 1820 -1950
rect 1840 -1970 1860 -1950
rect 1880 -1970 1900 -1950
rect 1920 -1970 1940 -1950
rect 1960 -1970 1980 -1950
rect 2000 -1970 2020 -1950
rect 2040 -1970 2060 -1950
rect 2080 -1970 2100 -1950
rect 2120 -1970 2140 -1950
rect 2160 -1970 2180 -1950
rect 2200 -1970 2220 -1950
rect 2240 -1970 2260 -1950
rect 2280 -1970 2300 -1950
rect 2320 -1970 2340 -1950
rect 2360 -1970 2380 -1950
rect 2400 -1970 2420 -1950
rect 2440 -1970 2460 -1950
rect 2480 -1970 2500 -1950
rect 2520 -1970 2540 -1950
rect 2560 -1970 2590 -1950
rect 120 -2065 140 -2045
rect 160 -2065 180 -2045
rect 200 -2065 220 -2045
rect 240 -2065 260 -2045
rect 280 -2065 300 -2045
rect 320 -2065 340 -2045
rect 360 -2065 380 -2045
rect 400 -2065 420 -2045
rect 440 -2065 460 -2045
rect 480 -2065 500 -2045
rect 520 -2065 540 -2045
rect 560 -2065 580 -2045
rect 600 -2065 620 -2045
rect 640 -2065 660 -2045
rect 680 -2065 700 -2045
rect 720 -2065 740 -2045
rect 760 -2065 780 -2045
rect 800 -2065 820 -2045
rect 840 -2065 860 -2045
rect 880 -2065 900 -2045
rect 920 -2065 940 -2045
rect 960 -2065 980 -2045
rect 1000 -2065 1020 -2045
rect 1040 -2065 1060 -2045
rect 1080 -2065 1100 -2045
rect 1120 -2065 1140 -2045
rect 1160 -2065 1180 -2045
rect 1200 -2065 1220 -2045
rect 1240 -2065 1260 -2045
rect 1280 -2065 1300 -2045
rect 1320 -2065 1340 -2045
rect 1360 -2065 1380 -2045
rect 1400 -2065 1420 -2045
rect 1440 -2065 1460 -2045
rect 1480 -2065 1500 -2045
rect 1520 -2065 1540 -2045
rect 1560 -2065 1580 -2045
rect 1600 -2065 1620 -2045
rect 1640 -2065 1660 -2045
rect 1680 -2065 1700 -2045
rect 1720 -2065 1740 -2045
rect 1760 -2065 1780 -2045
rect 1800 -2065 1820 -2045
rect 1840 -2065 1860 -2045
rect 1880 -2065 1900 -2045
rect 1920 -2065 1940 -2045
rect 1960 -2065 1980 -2045
rect 2000 -2065 2020 -2045
rect 2040 -2065 2060 -2045
rect 2080 -2065 2100 -2045
rect 2120 -2065 2140 -2045
rect 2160 -2065 2180 -2045
rect 2200 -2065 2220 -2045
rect 2240 -2065 2260 -2045
rect 2280 -2065 2300 -2045
rect 2320 -2065 2340 -2045
rect 2360 -2065 2380 -2045
rect 2400 -2065 2420 -2045
rect 2440 -2065 2460 -2045
rect 2480 -2065 2500 -2045
rect 2520 -2065 2540 -2045
rect 2560 -2065 2590 -2045
rect 120 -2160 140 -2140
rect 160 -2160 180 -2140
rect 200 -2160 220 -2140
rect 240 -2160 260 -2140
rect 280 -2160 300 -2140
rect 320 -2160 340 -2140
rect 360 -2160 380 -2140
rect 400 -2160 420 -2140
rect 440 -2160 460 -2140
rect 480 -2160 500 -2140
rect 520 -2160 540 -2140
rect 560 -2160 580 -2140
rect 600 -2160 620 -2140
rect 640 -2160 660 -2140
rect 680 -2160 700 -2140
rect 720 -2160 740 -2140
rect 760 -2160 780 -2140
rect 800 -2160 820 -2140
rect 840 -2160 860 -2140
rect 880 -2160 900 -2140
rect 920 -2160 940 -2140
rect 960 -2160 980 -2140
rect 1000 -2160 1020 -2140
rect 1040 -2160 1060 -2140
rect 1080 -2160 1100 -2140
rect 1120 -2160 1140 -2140
rect 1160 -2160 1180 -2140
rect 1200 -2160 1220 -2140
rect 1240 -2160 1260 -2140
rect 1280 -2160 1300 -2140
rect 1320 -2160 1340 -2140
rect 1360 -2160 1380 -2140
rect 1400 -2160 1420 -2140
rect 1440 -2160 1460 -2140
rect 1480 -2160 1500 -2140
rect 1520 -2160 1540 -2140
rect 1560 -2160 1580 -2140
rect 1600 -2160 1620 -2140
rect 1640 -2160 1660 -2140
rect 1680 -2160 1700 -2140
rect 1720 -2160 1740 -2140
rect 1760 -2160 1780 -2140
rect 1800 -2160 1820 -2140
rect 1840 -2160 1860 -2140
rect 1880 -2160 1900 -2140
rect 1920 -2160 1940 -2140
rect 1960 -2160 1980 -2140
rect 2000 -2160 2020 -2140
rect 2040 -2160 2060 -2140
rect 2080 -2160 2100 -2140
rect 2120 -2160 2140 -2140
rect 2160 -2160 2180 -2140
rect 2200 -2160 2220 -2140
rect 2240 -2160 2260 -2140
rect 2280 -2160 2300 -2140
rect 2320 -2160 2340 -2140
rect 2360 -2160 2380 -2140
rect 2400 -2160 2420 -2140
rect 2440 -2160 2460 -2140
rect 2480 -2160 2500 -2140
rect 2520 -2160 2540 -2140
rect 2560 -2160 2590 -2140
rect 120 -2255 140 -2235
rect 160 -2255 180 -2235
rect 200 -2255 220 -2235
rect 240 -2255 260 -2235
rect 280 -2255 300 -2235
rect 320 -2255 340 -2235
rect 360 -2255 380 -2235
rect 400 -2255 420 -2235
rect 440 -2255 460 -2235
rect 480 -2255 500 -2235
rect 520 -2255 540 -2235
rect 560 -2255 580 -2235
rect 600 -2255 620 -2235
rect 640 -2255 660 -2235
rect 680 -2255 700 -2235
rect 720 -2255 740 -2235
rect 760 -2255 780 -2235
rect 800 -2255 820 -2235
rect 840 -2255 860 -2235
rect 880 -2255 900 -2235
rect 920 -2255 940 -2235
rect 960 -2255 980 -2235
rect 1000 -2255 1020 -2235
rect 1040 -2255 1060 -2235
rect 1080 -2255 1100 -2235
rect 1120 -2255 1140 -2235
rect 1160 -2255 1180 -2235
rect 1200 -2255 1220 -2235
rect 1240 -2255 1260 -2235
rect 1280 -2255 1300 -2235
rect 1320 -2255 1340 -2235
rect 1360 -2255 1380 -2235
rect 1400 -2255 1420 -2235
rect 1440 -2255 1460 -2235
rect 1480 -2255 1500 -2235
rect 1520 -2255 1540 -2235
rect 1560 -2255 1580 -2235
rect 1600 -2255 1620 -2235
rect 1640 -2255 1660 -2235
rect 1680 -2255 1700 -2235
rect 1720 -2255 1740 -2235
rect 1760 -2255 1780 -2235
rect 1800 -2255 1820 -2235
rect 1840 -2255 1860 -2235
rect 1880 -2255 1900 -2235
rect 1920 -2255 1940 -2235
rect 1960 -2255 1980 -2235
rect 2000 -2255 2020 -2235
rect 2040 -2255 2060 -2235
rect 2080 -2255 2100 -2235
rect 2120 -2255 2140 -2235
rect 2160 -2255 2180 -2235
rect 2200 -2255 2220 -2235
rect 2240 -2255 2260 -2235
rect 2280 -2255 2300 -2235
rect 2320 -2255 2340 -2235
rect 2360 -2255 2380 -2235
rect 2400 -2255 2420 -2235
rect 2440 -2255 2460 -2235
rect 2480 -2255 2500 -2235
rect 2520 -2255 2540 -2235
rect 2560 -2255 2590 -2235
rect 120 -2350 140 -2330
rect 160 -2350 180 -2330
rect 200 -2350 220 -2330
rect 240 -2350 260 -2330
rect 280 -2350 300 -2330
rect 320 -2350 340 -2330
rect 360 -2350 380 -2330
rect 400 -2350 420 -2330
rect 440 -2350 460 -2330
rect 480 -2350 500 -2330
rect 520 -2350 540 -2330
rect 560 -2350 580 -2330
rect 600 -2350 620 -2330
rect 640 -2350 660 -2330
rect 680 -2350 700 -2330
rect 720 -2350 740 -2330
rect 760 -2350 780 -2330
rect 800 -2350 820 -2330
rect 840 -2350 860 -2330
rect 880 -2350 900 -2330
rect 920 -2350 940 -2330
rect 960 -2350 980 -2330
rect 1000 -2350 1020 -2330
rect 1040 -2350 1060 -2330
rect 1080 -2350 1100 -2330
rect 1120 -2350 1140 -2330
rect 1160 -2350 1180 -2330
rect 1200 -2350 1220 -2330
rect 1240 -2350 1260 -2330
rect 1280 -2350 1300 -2330
rect 1320 -2350 1340 -2330
rect 1360 -2350 1380 -2330
rect 1400 -2350 1420 -2330
rect 1440 -2350 1460 -2330
rect 1480 -2350 1500 -2330
rect 1520 -2350 1540 -2330
rect 1560 -2350 1580 -2330
rect 1600 -2350 1620 -2330
rect 1640 -2350 1660 -2330
rect 1680 -2350 1700 -2330
rect 1720 -2350 1740 -2330
rect 1760 -2350 1780 -2330
rect 1800 -2350 1820 -2330
rect 1840 -2350 1860 -2330
rect 1880 -2350 1900 -2330
rect 1920 -2350 1940 -2330
rect 1960 -2350 1980 -2330
rect 2000 -2350 2020 -2330
rect 2040 -2350 2060 -2330
rect 2080 -2350 2100 -2330
rect 2120 -2350 2140 -2330
rect 2160 -2350 2180 -2330
rect 2200 -2350 2220 -2330
rect 2240 -2350 2260 -2330
rect 2280 -2350 2300 -2330
rect 2320 -2350 2340 -2330
rect 2360 -2350 2380 -2330
rect 2400 -2350 2420 -2330
rect 2440 -2350 2460 -2330
rect 2480 -2350 2500 -2330
rect 2520 -2350 2540 -2330
rect 2560 -2350 2590 -2330
rect 120 -2445 140 -2425
rect 160 -2445 180 -2425
rect 200 -2445 220 -2425
rect 240 -2445 260 -2425
rect 280 -2445 300 -2425
rect 320 -2445 340 -2425
rect 360 -2445 380 -2425
rect 400 -2445 420 -2425
rect 440 -2445 460 -2425
rect 480 -2445 500 -2425
rect 520 -2445 540 -2425
rect 560 -2445 580 -2425
rect 600 -2445 620 -2425
rect 640 -2445 660 -2425
rect 680 -2445 700 -2425
rect 720 -2445 740 -2425
rect 760 -2445 780 -2425
rect 800 -2445 820 -2425
rect 840 -2445 860 -2425
rect 880 -2445 900 -2425
rect 920 -2445 940 -2425
rect 960 -2445 980 -2425
rect 1000 -2445 1020 -2425
rect 1040 -2445 1060 -2425
rect 1080 -2445 1100 -2425
rect 1120 -2445 1140 -2425
rect 1160 -2445 1180 -2425
rect 1200 -2445 1220 -2425
rect 1240 -2445 1260 -2425
rect 1280 -2445 1300 -2425
rect 1320 -2445 1340 -2425
rect 1360 -2445 1380 -2425
rect 1400 -2445 1420 -2425
rect 1440 -2445 1460 -2425
rect 1480 -2445 1500 -2425
rect 1520 -2445 1540 -2425
rect 1560 -2445 1580 -2425
rect 1600 -2445 1620 -2425
rect 1640 -2445 1660 -2425
rect 1680 -2445 1700 -2425
rect 1720 -2445 1740 -2425
rect 1760 -2445 1780 -2425
rect 1800 -2445 1820 -2425
rect 1840 -2445 1860 -2425
rect 1880 -2445 1900 -2425
rect 1920 -2445 1940 -2425
rect 1960 -2445 1980 -2425
rect 2000 -2445 2020 -2425
rect 2040 -2445 2060 -2425
rect 2080 -2445 2100 -2425
rect 2120 -2445 2140 -2425
rect 2160 -2445 2180 -2425
rect 2200 -2445 2220 -2425
rect 2240 -2445 2260 -2425
rect 2280 -2445 2300 -2425
rect 2320 -2445 2340 -2425
rect 2360 -2445 2380 -2425
rect 2400 -2445 2420 -2425
rect 2440 -2445 2460 -2425
rect 2480 -2445 2500 -2425
rect 2520 -2445 2540 -2425
rect 2560 -2445 2590 -2425
rect 120 -2540 140 -2520
rect 160 -2540 180 -2520
rect 200 -2540 220 -2520
rect 240 -2540 260 -2520
rect 280 -2540 300 -2520
rect 320 -2540 340 -2520
rect 360 -2540 380 -2520
rect 400 -2540 420 -2520
rect 440 -2540 460 -2520
rect 480 -2540 500 -2520
rect 520 -2540 540 -2520
rect 560 -2540 580 -2520
rect 600 -2540 620 -2520
rect 640 -2540 660 -2520
rect 680 -2540 700 -2520
rect 720 -2540 740 -2520
rect 760 -2540 780 -2520
rect 800 -2540 820 -2520
rect 840 -2540 860 -2520
rect 880 -2540 900 -2520
rect 920 -2540 940 -2520
rect 960 -2540 980 -2520
rect 1000 -2540 1020 -2520
rect 1040 -2540 1060 -2520
rect 1080 -2540 1100 -2520
rect 1120 -2540 1140 -2520
rect 1160 -2540 1180 -2520
rect 1200 -2540 1220 -2520
rect 1240 -2540 1260 -2520
rect 1280 -2540 1300 -2520
rect 1320 -2540 1340 -2520
rect 1360 -2540 1380 -2520
rect 1400 -2540 1420 -2520
rect 1440 -2540 1460 -2520
rect 1480 -2540 1500 -2520
rect 1520 -2540 1540 -2520
rect 1560 -2540 1580 -2520
rect 1600 -2540 1620 -2520
rect 1640 -2540 1660 -2520
rect 1680 -2540 1700 -2520
rect 1720 -2540 1740 -2520
rect 1760 -2540 1780 -2520
rect 1800 -2540 1820 -2520
rect 1840 -2540 1860 -2520
rect 1880 -2540 1900 -2520
rect 1920 -2540 1940 -2520
rect 1960 -2540 1980 -2520
rect 2000 -2540 2020 -2520
rect 2040 -2540 2060 -2520
rect 2080 -2540 2100 -2520
rect 2120 -2540 2140 -2520
rect 2160 -2540 2180 -2520
rect 2200 -2540 2220 -2520
rect 2240 -2540 2260 -2520
rect 2280 -2540 2300 -2520
rect 2320 -2540 2340 -2520
rect 2360 -2540 2380 -2520
rect 2400 -2540 2420 -2520
rect 2440 -2540 2460 -2520
rect 2480 -2540 2500 -2520
rect 2520 -2540 2540 -2520
rect 2560 -2540 2590 -2520
<< psubdiff >>
rect 175 2365 2675 2375
rect 175 2345 200 2365
rect 220 2345 240 2365
rect 260 2345 280 2365
rect 300 2345 320 2365
rect 340 2345 360 2365
rect 380 2345 400 2365
rect 420 2345 440 2365
rect 460 2345 480 2365
rect 500 2345 520 2365
rect 540 2345 560 2365
rect 580 2345 600 2365
rect 620 2345 640 2365
rect 660 2345 680 2365
rect 700 2345 720 2365
rect 740 2345 760 2365
rect 780 2345 800 2365
rect 820 2345 840 2365
rect 860 2345 880 2365
rect 900 2345 920 2365
rect 940 2345 960 2365
rect 980 2345 1000 2365
rect 1020 2345 1040 2365
rect 1060 2345 1080 2365
rect 1100 2345 1120 2365
rect 1140 2345 1160 2365
rect 1180 2345 1200 2365
rect 1220 2345 1240 2365
rect 1260 2345 1280 2365
rect 1300 2345 1320 2365
rect 1340 2345 1360 2365
rect 1380 2345 1400 2365
rect 1420 2345 1440 2365
rect 1460 2345 1480 2365
rect 1500 2345 1520 2365
rect 1540 2345 1560 2365
rect 1580 2345 1600 2365
rect 1620 2345 1640 2365
rect 1660 2345 1680 2365
rect 1700 2345 1720 2365
rect 1740 2345 1760 2365
rect 1780 2345 1800 2365
rect 1820 2345 1840 2365
rect 1860 2345 1880 2365
rect 1900 2345 1920 2365
rect 1940 2345 1960 2365
rect 1980 2345 2000 2365
rect 2020 2345 2040 2365
rect 2060 2345 2080 2365
rect 2100 2345 2120 2365
rect 2140 2345 2160 2365
rect 2180 2345 2200 2365
rect 2220 2345 2240 2365
rect 2260 2345 2280 2365
rect 2300 2345 2320 2365
rect 2340 2345 2360 2365
rect 2380 2345 2400 2365
rect 2420 2345 2440 2365
rect 2460 2345 2480 2365
rect 2500 2345 2520 2365
rect 2540 2345 2560 2365
rect 2580 2345 2600 2365
rect 2620 2345 2640 2365
rect 2660 2345 2675 2365
rect 175 2335 2675 2345
rect 175 95 2675 105
rect 175 75 200 95
rect 220 75 240 95
rect 260 75 280 95
rect 300 75 320 95
rect 340 75 360 95
rect 380 75 400 95
rect 420 75 440 95
rect 460 75 480 95
rect 500 75 520 95
rect 540 75 560 95
rect 580 75 600 95
rect 620 75 640 95
rect 660 75 680 95
rect 700 75 720 95
rect 740 75 760 95
rect 780 75 800 95
rect 820 75 840 95
rect 860 75 880 95
rect 900 75 920 95
rect 940 75 960 95
rect 980 75 1000 95
rect 1020 75 1040 95
rect 1060 75 1080 95
rect 1100 75 1120 95
rect 1140 75 1160 95
rect 1180 75 1200 95
rect 1220 75 1240 95
rect 1260 75 1280 95
rect 1300 75 1320 95
rect 1340 75 1360 95
rect 1380 75 1400 95
rect 1420 75 1440 95
rect 1460 75 1480 95
rect 1500 75 1520 95
rect 1540 75 1560 95
rect 1580 75 1600 95
rect 1620 75 1640 95
rect 1660 75 1680 95
rect 1700 75 1720 95
rect 1740 75 1760 95
rect 1780 75 1800 95
rect 1820 75 1840 95
rect 1860 75 1880 95
rect 1900 75 1920 95
rect 1940 75 1960 95
rect 1980 75 2000 95
rect 2020 75 2040 95
rect 2060 75 2080 95
rect 2100 75 2120 95
rect 2140 75 2160 95
rect 2180 75 2200 95
rect 2220 75 2240 95
rect 2260 75 2280 95
rect 2300 75 2320 95
rect 2340 75 2360 95
rect 2380 75 2400 95
rect 2420 75 2440 95
rect 2460 75 2480 95
rect 2500 75 2520 95
rect 2540 75 2560 95
rect 2580 75 2600 95
rect 2620 75 2640 95
rect 2660 75 2675 95
rect 175 65 2675 75
rect 105 -10 2605 0
rect 105 -30 120 -10
rect 140 -30 160 -10
rect 180 -30 200 -10
rect 220 -30 240 -10
rect 260 -30 280 -10
rect 300 -30 320 -10
rect 340 -30 360 -10
rect 380 -30 400 -10
rect 420 -30 440 -10
rect 460 -30 480 -10
rect 500 -30 520 -10
rect 540 -30 560 -10
rect 580 -30 600 -10
rect 620 -30 640 -10
rect 660 -30 680 -10
rect 700 -30 720 -10
rect 740 -30 760 -10
rect 780 -30 800 -10
rect 820 -30 840 -10
rect 860 -30 880 -10
rect 900 -30 920 -10
rect 940 -30 960 -10
rect 980 -30 1000 -10
rect 1020 -30 1040 -10
rect 1060 -30 1080 -10
rect 1100 -30 1120 -10
rect 1140 -30 1160 -10
rect 1180 -30 1200 -10
rect 1220 -30 1240 -10
rect 1260 -30 1280 -10
rect 1300 -30 1320 -10
rect 1340 -30 1360 -10
rect 1380 -30 1400 -10
rect 1420 -30 1440 -10
rect 1460 -30 1480 -10
rect 1500 -30 1520 -10
rect 1540 -30 1560 -10
rect 1580 -30 1600 -10
rect 1620 -30 1640 -10
rect 1660 -30 1680 -10
rect 1700 -30 1720 -10
rect 1740 -30 1760 -10
rect 1780 -30 1800 -10
rect 1820 -30 1840 -10
rect 1860 -30 1880 -10
rect 1900 -30 1920 -10
rect 1940 -30 1960 -10
rect 1980 -30 2000 -10
rect 2020 -30 2040 -10
rect 2060 -30 2080 -10
rect 2100 -30 2120 -10
rect 2140 -30 2160 -10
rect 2180 -30 2200 -10
rect 2220 -30 2240 -10
rect 2260 -30 2280 -10
rect 2300 -30 2320 -10
rect 2340 -30 2360 -10
rect 2380 -30 2400 -10
rect 2420 -30 2440 -10
rect 2460 -30 2480 -10
rect 2500 -30 2520 -10
rect 2540 -30 2560 -10
rect 2590 -30 2605 -10
rect 105 -40 2605 -30
rect 105 -2560 2605 -2550
rect 105 -2580 120 -2560
rect 140 -2580 160 -2560
rect 180 -2580 200 -2560
rect 220 -2580 240 -2560
rect 260 -2580 280 -2560
rect 300 -2580 320 -2560
rect 340 -2580 360 -2560
rect 380 -2580 400 -2560
rect 420 -2580 440 -2560
rect 460 -2580 480 -2560
rect 500 -2580 520 -2560
rect 540 -2580 560 -2560
rect 580 -2580 600 -2560
rect 620 -2580 640 -2560
rect 660 -2580 680 -2560
rect 700 -2580 720 -2560
rect 740 -2580 760 -2560
rect 780 -2580 800 -2560
rect 820 -2580 840 -2560
rect 860 -2580 880 -2560
rect 900 -2580 920 -2560
rect 940 -2580 960 -2560
rect 980 -2580 1000 -2560
rect 1020 -2580 1040 -2560
rect 1060 -2580 1080 -2560
rect 1100 -2580 1120 -2560
rect 1140 -2580 1160 -2560
rect 1180 -2580 1200 -2560
rect 1220 -2580 1240 -2560
rect 1260 -2580 1280 -2560
rect 1300 -2580 1320 -2560
rect 1340 -2580 1360 -2560
rect 1380 -2580 1400 -2560
rect 1420 -2580 1440 -2560
rect 1460 -2580 1480 -2560
rect 1500 -2580 1520 -2560
rect 1540 -2580 1560 -2560
rect 1580 -2580 1600 -2560
rect 1620 -2580 1640 -2560
rect 1660 -2580 1680 -2560
rect 1700 -2580 1720 -2560
rect 1740 -2580 1760 -2560
rect 1780 -2580 1800 -2560
rect 1820 -2580 1840 -2560
rect 1860 -2580 1880 -2560
rect 1900 -2580 1920 -2560
rect 1940 -2580 1960 -2560
rect 1980 -2580 2000 -2560
rect 2020 -2580 2040 -2560
rect 2060 -2580 2080 -2560
rect 2100 -2580 2120 -2560
rect 2140 -2580 2160 -2560
rect 2180 -2580 2200 -2560
rect 2220 -2580 2240 -2560
rect 2260 -2580 2280 -2560
rect 2300 -2580 2320 -2560
rect 2340 -2580 2360 -2560
rect 2380 -2580 2400 -2560
rect 2420 -2580 2440 -2560
rect 2460 -2580 2480 -2560
rect 2500 -2580 2520 -2560
rect 2540 -2580 2560 -2560
rect 2590 -2580 2605 -2560
rect 105 -2590 2605 -2580
<< psubdiffcont >>
rect 200 2345 220 2365
rect 240 2345 260 2365
rect 280 2345 300 2365
rect 320 2345 340 2365
rect 360 2345 380 2365
rect 400 2345 420 2365
rect 440 2345 460 2365
rect 480 2345 500 2365
rect 520 2345 540 2365
rect 560 2345 580 2365
rect 600 2345 620 2365
rect 640 2345 660 2365
rect 680 2345 700 2365
rect 720 2345 740 2365
rect 760 2345 780 2365
rect 800 2345 820 2365
rect 840 2345 860 2365
rect 880 2345 900 2365
rect 920 2345 940 2365
rect 960 2345 980 2365
rect 1000 2345 1020 2365
rect 1040 2345 1060 2365
rect 1080 2345 1100 2365
rect 1120 2345 1140 2365
rect 1160 2345 1180 2365
rect 1200 2345 1220 2365
rect 1240 2345 1260 2365
rect 1280 2345 1300 2365
rect 1320 2345 1340 2365
rect 1360 2345 1380 2365
rect 1400 2345 1420 2365
rect 1440 2345 1460 2365
rect 1480 2345 1500 2365
rect 1520 2345 1540 2365
rect 1560 2345 1580 2365
rect 1600 2345 1620 2365
rect 1640 2345 1660 2365
rect 1680 2345 1700 2365
rect 1720 2345 1740 2365
rect 1760 2345 1780 2365
rect 1800 2345 1820 2365
rect 1840 2345 1860 2365
rect 1880 2345 1900 2365
rect 1920 2345 1940 2365
rect 1960 2345 1980 2365
rect 2000 2345 2020 2365
rect 2040 2345 2060 2365
rect 2080 2345 2100 2365
rect 2120 2345 2140 2365
rect 2160 2345 2180 2365
rect 2200 2345 2220 2365
rect 2240 2345 2260 2365
rect 2280 2345 2300 2365
rect 2320 2345 2340 2365
rect 2360 2345 2380 2365
rect 2400 2345 2420 2365
rect 2440 2345 2460 2365
rect 2480 2345 2500 2365
rect 2520 2345 2540 2365
rect 2560 2345 2580 2365
rect 2600 2345 2620 2365
rect 2640 2345 2660 2365
rect 200 75 220 95
rect 240 75 260 95
rect 280 75 300 95
rect 320 75 340 95
rect 360 75 380 95
rect 400 75 420 95
rect 440 75 460 95
rect 480 75 500 95
rect 520 75 540 95
rect 560 75 580 95
rect 600 75 620 95
rect 640 75 660 95
rect 680 75 700 95
rect 720 75 740 95
rect 760 75 780 95
rect 800 75 820 95
rect 840 75 860 95
rect 880 75 900 95
rect 920 75 940 95
rect 960 75 980 95
rect 1000 75 1020 95
rect 1040 75 1060 95
rect 1080 75 1100 95
rect 1120 75 1140 95
rect 1160 75 1180 95
rect 1200 75 1220 95
rect 1240 75 1260 95
rect 1280 75 1300 95
rect 1320 75 1340 95
rect 1360 75 1380 95
rect 1400 75 1420 95
rect 1440 75 1460 95
rect 1480 75 1500 95
rect 1520 75 1540 95
rect 1560 75 1580 95
rect 1600 75 1620 95
rect 1640 75 1660 95
rect 1680 75 1700 95
rect 1720 75 1740 95
rect 1760 75 1780 95
rect 1800 75 1820 95
rect 1840 75 1860 95
rect 1880 75 1900 95
rect 1920 75 1940 95
rect 1960 75 1980 95
rect 2000 75 2020 95
rect 2040 75 2060 95
rect 2080 75 2100 95
rect 2120 75 2140 95
rect 2160 75 2180 95
rect 2200 75 2220 95
rect 2240 75 2260 95
rect 2280 75 2300 95
rect 2320 75 2340 95
rect 2360 75 2380 95
rect 2400 75 2420 95
rect 2440 75 2460 95
rect 2480 75 2500 95
rect 2520 75 2540 95
rect 2560 75 2580 95
rect 2600 75 2620 95
rect 2640 75 2660 95
rect 120 -30 140 -10
rect 160 -30 180 -10
rect 200 -30 220 -10
rect 240 -30 260 -10
rect 280 -30 300 -10
rect 320 -30 340 -10
rect 360 -30 380 -10
rect 400 -30 420 -10
rect 440 -30 460 -10
rect 480 -30 500 -10
rect 520 -30 540 -10
rect 560 -30 580 -10
rect 600 -30 620 -10
rect 640 -30 660 -10
rect 680 -30 700 -10
rect 720 -30 740 -10
rect 760 -30 780 -10
rect 800 -30 820 -10
rect 840 -30 860 -10
rect 880 -30 900 -10
rect 920 -30 940 -10
rect 960 -30 980 -10
rect 1000 -30 1020 -10
rect 1040 -30 1060 -10
rect 1080 -30 1100 -10
rect 1120 -30 1140 -10
rect 1160 -30 1180 -10
rect 1200 -30 1220 -10
rect 1240 -30 1260 -10
rect 1280 -30 1300 -10
rect 1320 -30 1340 -10
rect 1360 -30 1380 -10
rect 1400 -30 1420 -10
rect 1440 -30 1460 -10
rect 1480 -30 1500 -10
rect 1520 -30 1540 -10
rect 1560 -30 1580 -10
rect 1600 -30 1620 -10
rect 1640 -30 1660 -10
rect 1680 -30 1700 -10
rect 1720 -30 1740 -10
rect 1760 -30 1780 -10
rect 1800 -30 1820 -10
rect 1840 -30 1860 -10
rect 1880 -30 1900 -10
rect 1920 -30 1940 -10
rect 1960 -30 1980 -10
rect 2000 -30 2020 -10
rect 2040 -30 2060 -10
rect 2080 -30 2100 -10
rect 2120 -30 2140 -10
rect 2160 -30 2180 -10
rect 2200 -30 2220 -10
rect 2240 -30 2260 -10
rect 2280 -30 2300 -10
rect 2320 -30 2340 -10
rect 2360 -30 2380 -10
rect 2400 -30 2420 -10
rect 2440 -30 2460 -10
rect 2480 -30 2500 -10
rect 2520 -30 2540 -10
rect 2560 -30 2590 -10
rect 120 -2580 140 -2560
rect 160 -2580 180 -2560
rect 200 -2580 220 -2560
rect 240 -2580 260 -2560
rect 280 -2580 300 -2560
rect 320 -2580 340 -2560
rect 360 -2580 380 -2560
rect 400 -2580 420 -2560
rect 440 -2580 460 -2560
rect 480 -2580 500 -2560
rect 520 -2580 540 -2560
rect 560 -2580 580 -2560
rect 600 -2580 620 -2560
rect 640 -2580 660 -2560
rect 680 -2580 700 -2560
rect 720 -2580 740 -2560
rect 760 -2580 780 -2560
rect 800 -2580 820 -2560
rect 840 -2580 860 -2560
rect 880 -2580 900 -2560
rect 920 -2580 940 -2560
rect 960 -2580 980 -2560
rect 1000 -2580 1020 -2560
rect 1040 -2580 1060 -2560
rect 1080 -2580 1100 -2560
rect 1120 -2580 1140 -2560
rect 1160 -2580 1180 -2560
rect 1200 -2580 1220 -2560
rect 1240 -2580 1260 -2560
rect 1280 -2580 1300 -2560
rect 1320 -2580 1340 -2560
rect 1360 -2580 1380 -2560
rect 1400 -2580 1420 -2560
rect 1440 -2580 1460 -2560
rect 1480 -2580 1500 -2560
rect 1520 -2580 1540 -2560
rect 1560 -2580 1580 -2560
rect 1600 -2580 1620 -2560
rect 1640 -2580 1660 -2560
rect 1680 -2580 1700 -2560
rect 1720 -2580 1740 -2560
rect 1760 -2580 1780 -2560
rect 1800 -2580 1820 -2560
rect 1840 -2580 1860 -2560
rect 1880 -2580 1900 -2560
rect 1920 -2580 1940 -2560
rect 1960 -2580 1980 -2560
rect 2000 -2580 2020 -2560
rect 2040 -2580 2060 -2560
rect 2080 -2580 2100 -2560
rect 2120 -2580 2140 -2560
rect 2160 -2580 2180 -2560
rect 2200 -2580 2220 -2560
rect 2240 -2580 2260 -2560
rect 2280 -2580 2300 -2560
rect 2320 -2580 2340 -2560
rect 2360 -2580 2380 -2560
rect 2400 -2580 2420 -2560
rect 2440 -2580 2460 -2560
rect 2480 -2580 2500 -2560
rect 2520 -2580 2540 -2560
rect 2560 -2580 2590 -2560
<< poly >>
rect 0 2262 165 2265
rect 0 2255 175 2262
rect 0 2235 10 2255
rect 30 2235 50 2255
rect 70 2235 90 2255
rect 110 2235 130 2255
rect 155 2235 175 2255
rect 0 2230 175 2235
rect 2675 2230 2690 2262
rect 0 2225 165 2230
rect 0 2180 165 2185
rect 0 2175 175 2180
rect 0 2155 10 2175
rect 30 2155 50 2175
rect 70 2155 90 2175
rect 110 2155 130 2175
rect 155 2155 175 2175
rect 0 2148 175 2155
rect 2675 2148 2690 2180
rect 0 2145 165 2148
rect 0 2098 165 2100
rect 0 2090 175 2098
rect 0 2070 10 2090
rect 30 2070 50 2090
rect 70 2070 90 2090
rect 110 2070 130 2090
rect 155 2070 175 2090
rect 0 2066 175 2070
rect 2675 2066 2690 2098
rect 0 2060 165 2066
rect 0 2016 165 2020
rect 0 2010 175 2016
rect 0 1990 10 2010
rect 30 1990 50 2010
rect 70 1990 90 2010
rect 110 1990 130 2010
rect 155 1990 175 2010
rect 0 1984 175 1990
rect 2675 1984 2690 2016
rect 0 1980 165 1984
rect 0 1934 165 1940
rect 0 1930 175 1934
rect 0 1910 10 1930
rect 30 1910 50 1930
rect 70 1910 90 1930
rect 110 1910 130 1930
rect 155 1910 175 1930
rect 0 1902 175 1910
rect 2675 1902 2690 1934
rect 0 1900 165 1902
rect 0 1852 165 1855
rect 0 1845 175 1852
rect 0 1825 10 1845
rect 30 1825 50 1845
rect 70 1825 90 1845
rect 110 1825 130 1845
rect 155 1825 175 1845
rect 0 1820 175 1825
rect 2675 1820 2690 1852
rect 0 1815 165 1820
rect 0 1770 165 1775
rect 0 1765 175 1770
rect 0 1745 10 1765
rect 30 1745 50 1765
rect 70 1745 90 1765
rect 110 1745 130 1765
rect 155 1745 175 1765
rect 0 1738 175 1745
rect 2675 1738 2690 1770
rect 0 1735 165 1738
rect 0 1688 165 1690
rect 0 1680 175 1688
rect 0 1660 10 1680
rect 30 1660 50 1680
rect 70 1660 90 1680
rect 110 1660 130 1680
rect 155 1660 175 1680
rect 0 1656 175 1660
rect 2675 1656 2690 1688
rect 0 1650 165 1656
rect 0 1606 165 1610
rect 0 1600 175 1606
rect 0 1580 10 1600
rect 30 1580 50 1600
rect 70 1580 90 1600
rect 110 1580 130 1600
rect 155 1580 175 1600
rect 0 1574 175 1580
rect 2675 1574 2690 1606
rect 0 1570 165 1574
rect 0 1524 165 1530
rect 0 1520 175 1524
rect 0 1500 10 1520
rect 30 1500 50 1520
rect 70 1500 90 1520
rect 110 1500 130 1520
rect 155 1500 175 1520
rect 0 1492 175 1500
rect 2675 1492 2690 1524
rect 0 1490 165 1492
rect 0 1442 165 1445
rect 0 1435 175 1442
rect 0 1415 10 1435
rect 30 1415 50 1435
rect 70 1415 90 1435
rect 110 1415 130 1435
rect 155 1415 175 1435
rect 0 1410 175 1415
rect 2675 1410 2690 1442
rect 0 1405 165 1410
rect 0 1360 165 1365
rect 0 1355 175 1360
rect 0 1335 10 1355
rect 30 1335 50 1355
rect 70 1335 90 1355
rect 110 1335 130 1355
rect 155 1335 175 1355
rect 0 1328 175 1335
rect 2675 1328 2690 1360
rect 0 1325 165 1328
rect 0 1278 165 1280
rect 0 1270 175 1278
rect 0 1250 10 1270
rect 30 1250 50 1270
rect 70 1250 90 1270
rect 110 1250 130 1270
rect 155 1250 175 1270
rect 0 1246 175 1250
rect 2675 1246 2690 1278
rect 0 1240 165 1246
rect 0 1196 165 1200
rect 0 1190 175 1196
rect 0 1170 10 1190
rect 30 1170 50 1190
rect 70 1170 90 1190
rect 110 1170 130 1190
rect 155 1170 175 1190
rect 0 1164 175 1170
rect 2675 1164 2690 1196
rect 0 1160 165 1164
rect 0 1114 165 1120
rect 0 1110 175 1114
rect 0 1090 10 1110
rect 30 1090 50 1110
rect 70 1090 90 1110
rect 110 1090 130 1110
rect 155 1090 175 1110
rect 0 1082 175 1090
rect 2675 1082 2690 1114
rect 0 1080 165 1082
rect 0 1032 165 1035
rect 0 1025 175 1032
rect 0 1005 10 1025
rect 30 1005 50 1025
rect 70 1005 90 1025
rect 110 1005 130 1025
rect 155 1005 175 1025
rect 0 1000 175 1005
rect 2675 1000 2690 1032
rect 0 995 165 1000
rect 0 950 165 955
rect 0 945 175 950
rect 0 925 10 945
rect 30 925 50 945
rect 70 925 90 945
rect 110 925 130 945
rect 155 925 175 945
rect 0 918 175 925
rect 2675 918 2690 950
rect 0 915 165 918
rect 0 868 165 870
rect 0 860 175 868
rect 0 840 10 860
rect 30 840 50 860
rect 70 840 90 860
rect 110 840 130 860
rect 155 840 175 860
rect 0 836 175 840
rect 2675 836 2690 868
rect 0 830 165 836
rect 0 786 165 790
rect 0 780 175 786
rect 0 760 10 780
rect 30 760 50 780
rect 70 760 90 780
rect 110 760 130 780
rect 155 760 175 780
rect 0 754 175 760
rect 2675 754 2690 786
rect 0 750 165 754
rect 0 704 165 710
rect 0 700 175 704
rect 0 680 10 700
rect 30 680 50 700
rect 70 680 90 700
rect 110 680 130 700
rect 155 680 175 700
rect 0 672 175 680
rect 2675 672 2690 704
rect 0 670 165 672
rect 0 622 165 625
rect 0 615 175 622
rect 0 595 10 615
rect 30 595 50 615
rect 70 595 90 615
rect 110 595 130 615
rect 155 595 175 615
rect 0 590 175 595
rect 2675 590 2690 622
rect 0 585 165 590
rect 0 540 165 545
rect 0 535 175 540
rect 0 515 10 535
rect 30 515 50 535
rect 70 515 90 535
rect 110 515 130 535
rect 155 515 175 535
rect 0 508 175 515
rect 2675 508 2690 540
rect 0 505 165 508
rect 0 458 165 465
rect 0 455 175 458
rect 0 435 10 455
rect 30 435 50 455
rect 70 435 90 455
rect 110 435 130 455
rect 155 435 175 455
rect 0 426 175 435
rect 2675 426 2690 458
rect 0 425 165 426
rect 0 376 165 380
rect 0 370 175 376
rect 0 350 10 370
rect 30 350 50 370
rect 70 350 90 370
rect 110 350 130 370
rect 155 350 175 370
rect 0 344 175 350
rect 2675 344 2690 376
rect 0 340 165 344
rect 0 294 165 300
rect 0 290 175 294
rect 0 270 10 290
rect 30 270 50 290
rect 70 270 90 290
rect 110 270 130 290
rect 155 270 175 290
rect 0 262 175 270
rect 2675 262 2690 294
rect 0 260 165 262
rect 0 212 165 220
rect 0 210 175 212
rect 0 190 10 210
rect 30 190 50 210
rect 70 190 90 210
rect 110 190 130 210
rect 155 190 175 210
rect 0 180 175 190
rect 2675 180 2690 212
rect -70 -95 105 -85
rect -70 -120 -60 -95
rect -40 -120 -20 -95
rect 0 -120 20 -95
rect 40 -120 60 -95
rect 85 -120 105 -95
rect -70 -130 105 -120
rect 2605 -130 2620 -85
rect -70 -190 105 -180
rect -70 -215 -60 -190
rect -40 -215 -20 -190
rect 0 -215 20 -190
rect 40 -215 60 -190
rect 85 -215 105 -190
rect -70 -225 105 -215
rect 2605 -225 2620 -180
rect -70 -285 105 -275
rect -70 -310 -60 -285
rect -40 -310 -20 -285
rect 0 -310 20 -285
rect 40 -310 60 -285
rect 85 -310 105 -285
rect -70 -320 105 -310
rect 2605 -320 2620 -275
rect -70 -380 105 -370
rect -70 -405 -60 -380
rect -40 -405 -20 -380
rect 0 -405 20 -380
rect 40 -405 60 -380
rect 85 -405 105 -380
rect -70 -415 105 -405
rect 2605 -415 2620 -370
rect -70 -475 105 -465
rect -70 -500 -60 -475
rect -40 -500 -20 -475
rect 0 -500 20 -475
rect 40 -500 60 -475
rect 85 -500 105 -475
rect -70 -510 105 -500
rect 2605 -510 2620 -465
rect -70 -570 105 -560
rect -70 -595 -60 -570
rect -40 -595 -20 -570
rect 0 -595 20 -570
rect 40 -595 60 -570
rect 85 -595 105 -570
rect -70 -605 105 -595
rect 2605 -605 2620 -560
rect -70 -665 105 -655
rect -70 -690 -60 -665
rect -40 -690 -20 -665
rect 0 -690 20 -665
rect 40 -690 60 -665
rect 85 -690 105 -665
rect -70 -700 105 -690
rect 2605 -700 2620 -655
rect -70 -760 105 -750
rect -70 -785 -60 -760
rect -40 -785 -20 -760
rect 0 -785 20 -760
rect 40 -785 60 -760
rect 85 -785 105 -760
rect -70 -795 105 -785
rect 2605 -795 2620 -750
rect -70 -855 105 -845
rect -70 -880 -60 -855
rect -40 -880 -20 -855
rect 0 -880 20 -855
rect 40 -880 60 -855
rect 85 -880 105 -855
rect -70 -890 105 -880
rect 2605 -890 2620 -845
rect -70 -950 105 -940
rect -70 -975 -60 -950
rect -40 -975 -20 -950
rect 0 -975 20 -950
rect 40 -975 60 -950
rect 85 -975 105 -950
rect -70 -985 105 -975
rect 2605 -985 2620 -940
rect -70 -1045 105 -1035
rect -70 -1070 -60 -1045
rect -40 -1070 -20 -1045
rect 0 -1070 20 -1045
rect 40 -1070 60 -1045
rect 85 -1070 105 -1045
rect -70 -1080 105 -1070
rect 2605 -1080 2620 -1035
rect -70 -1140 105 -1130
rect -70 -1165 -60 -1140
rect -40 -1165 -20 -1140
rect 0 -1165 20 -1140
rect 40 -1165 60 -1140
rect 85 -1165 105 -1140
rect -70 -1175 105 -1165
rect 2605 -1175 2620 -1130
rect -70 -1235 105 -1225
rect -70 -1260 -60 -1235
rect -40 -1260 -20 -1235
rect 0 -1260 20 -1235
rect 40 -1260 60 -1235
rect 85 -1260 105 -1235
rect -70 -1270 105 -1260
rect 2605 -1270 2620 -1225
rect -70 -1330 105 -1320
rect -70 -1355 -60 -1330
rect -40 -1355 -20 -1330
rect 0 -1355 20 -1330
rect 40 -1355 60 -1330
rect 85 -1355 105 -1330
rect -70 -1365 105 -1355
rect 2605 -1365 2620 -1320
rect -70 -1425 105 -1415
rect -70 -1450 -60 -1425
rect -40 -1450 -20 -1425
rect 0 -1450 20 -1425
rect 40 -1450 60 -1425
rect 85 -1450 105 -1425
rect -70 -1460 105 -1450
rect 2605 -1460 2620 -1415
rect -70 -1520 105 -1510
rect -70 -1545 -60 -1520
rect -40 -1545 -20 -1520
rect 0 -1545 20 -1520
rect 40 -1545 60 -1520
rect 85 -1545 105 -1520
rect -70 -1555 105 -1545
rect 2605 -1555 2620 -1510
rect -70 -1615 105 -1605
rect -70 -1640 -60 -1615
rect -40 -1640 -20 -1615
rect 0 -1640 20 -1615
rect 40 -1640 60 -1615
rect 85 -1640 105 -1615
rect -70 -1650 105 -1640
rect 2605 -1650 2620 -1605
rect -70 -1710 105 -1700
rect -70 -1735 -60 -1710
rect -40 -1735 -20 -1710
rect 0 -1735 20 -1710
rect 40 -1735 60 -1710
rect 85 -1735 105 -1710
rect -70 -1745 105 -1735
rect 2605 -1745 2620 -1700
rect -70 -1805 105 -1795
rect -70 -1830 -60 -1805
rect -40 -1830 -20 -1805
rect 0 -1830 20 -1805
rect 40 -1830 60 -1805
rect 85 -1830 105 -1805
rect -70 -1840 105 -1830
rect 2605 -1840 2620 -1795
rect -70 -1900 105 -1890
rect -70 -1925 -60 -1900
rect -40 -1925 -20 -1900
rect 0 -1925 20 -1900
rect 40 -1925 60 -1900
rect 85 -1925 105 -1900
rect -70 -1935 105 -1925
rect 2605 -1935 2620 -1890
rect -70 -1995 105 -1985
rect -70 -2020 -60 -1995
rect -40 -2020 -20 -1995
rect 0 -2020 20 -1995
rect 40 -2020 60 -1995
rect 85 -2020 105 -1995
rect -70 -2030 105 -2020
rect 2605 -2030 2620 -1985
rect -70 -2090 105 -2080
rect -70 -2115 -60 -2090
rect -40 -2115 -20 -2090
rect 0 -2115 20 -2090
rect 40 -2115 60 -2090
rect 85 -2115 105 -2090
rect -70 -2125 105 -2115
rect 2605 -2125 2620 -2080
rect -70 -2185 105 -2175
rect -70 -2210 -60 -2185
rect -40 -2210 -20 -2185
rect 0 -2210 20 -2185
rect 40 -2210 60 -2185
rect 85 -2210 105 -2185
rect -70 -2220 105 -2210
rect 2605 -2220 2620 -2175
rect -70 -2280 105 -2270
rect -70 -2305 -60 -2280
rect -40 -2305 -20 -2280
rect 0 -2305 20 -2280
rect 40 -2305 60 -2280
rect 85 -2305 105 -2280
rect -70 -2315 105 -2305
rect 2605 -2315 2620 -2270
rect -70 -2375 105 -2365
rect -70 -2400 -60 -2375
rect -40 -2400 -20 -2375
rect 0 -2400 20 -2375
rect 40 -2400 60 -2375
rect 85 -2400 105 -2375
rect -70 -2410 105 -2400
rect 2605 -2410 2620 -2365
rect -70 -2470 105 -2460
rect -70 -2495 -60 -2470
rect -40 -2495 -20 -2470
rect 0 -2495 20 -2470
rect 40 -2495 60 -2470
rect 85 -2495 105 -2470
rect -70 -2505 105 -2495
rect 2605 -2505 2620 -2460
<< polycont >>
rect 10 2235 30 2255
rect 50 2235 70 2255
rect 90 2235 110 2255
rect 130 2235 155 2255
rect 10 2155 30 2175
rect 50 2155 70 2175
rect 90 2155 110 2175
rect 130 2155 155 2175
rect 10 2070 30 2090
rect 50 2070 70 2090
rect 90 2070 110 2090
rect 130 2070 155 2090
rect 10 1990 30 2010
rect 50 1990 70 2010
rect 90 1990 110 2010
rect 130 1990 155 2010
rect 10 1910 30 1930
rect 50 1910 70 1930
rect 90 1910 110 1930
rect 130 1910 155 1930
rect 10 1825 30 1845
rect 50 1825 70 1845
rect 90 1825 110 1845
rect 130 1825 155 1845
rect 10 1745 30 1765
rect 50 1745 70 1765
rect 90 1745 110 1765
rect 130 1745 155 1765
rect 10 1660 30 1680
rect 50 1660 70 1680
rect 90 1660 110 1680
rect 130 1660 155 1680
rect 10 1580 30 1600
rect 50 1580 70 1600
rect 90 1580 110 1600
rect 130 1580 155 1600
rect 10 1500 30 1520
rect 50 1500 70 1520
rect 90 1500 110 1520
rect 130 1500 155 1520
rect 10 1415 30 1435
rect 50 1415 70 1435
rect 90 1415 110 1435
rect 130 1415 155 1435
rect 10 1335 30 1355
rect 50 1335 70 1355
rect 90 1335 110 1355
rect 130 1335 155 1355
rect 10 1250 30 1270
rect 50 1250 70 1270
rect 90 1250 110 1270
rect 130 1250 155 1270
rect 10 1170 30 1190
rect 50 1170 70 1190
rect 90 1170 110 1190
rect 130 1170 155 1190
rect 10 1090 30 1110
rect 50 1090 70 1110
rect 90 1090 110 1110
rect 130 1090 155 1110
rect 10 1005 30 1025
rect 50 1005 70 1025
rect 90 1005 110 1025
rect 130 1005 155 1025
rect 10 925 30 945
rect 50 925 70 945
rect 90 925 110 945
rect 130 925 155 945
rect 10 840 30 860
rect 50 840 70 860
rect 90 840 110 860
rect 130 840 155 860
rect 10 760 30 780
rect 50 760 70 780
rect 90 760 110 780
rect 130 760 155 780
rect 10 680 30 700
rect 50 680 70 700
rect 90 680 110 700
rect 130 680 155 700
rect 10 595 30 615
rect 50 595 70 615
rect 90 595 110 615
rect 130 595 155 615
rect 10 515 30 535
rect 50 515 70 535
rect 90 515 110 535
rect 130 515 155 535
rect 10 435 30 455
rect 50 435 70 455
rect 90 435 110 455
rect 130 435 155 455
rect 10 350 30 370
rect 50 350 70 370
rect 90 350 110 370
rect 130 350 155 370
rect 10 270 30 290
rect 50 270 70 290
rect 90 270 110 290
rect 130 270 155 290
rect 10 190 30 210
rect 50 190 70 210
rect 90 190 110 210
rect 130 190 155 210
rect -60 -120 -40 -95
rect -20 -120 0 -95
rect 20 -120 40 -95
rect 60 -120 85 -95
rect -60 -215 -40 -190
rect -20 -215 0 -190
rect 20 -215 40 -190
rect 60 -215 85 -190
rect -60 -310 -40 -285
rect -20 -310 0 -285
rect 20 -310 40 -285
rect 60 -310 85 -285
rect -60 -405 -40 -380
rect -20 -405 0 -380
rect 20 -405 40 -380
rect 60 -405 85 -380
rect -60 -500 -40 -475
rect -20 -500 0 -475
rect 20 -500 40 -475
rect 60 -500 85 -475
rect -60 -595 -40 -570
rect -20 -595 0 -570
rect 20 -595 40 -570
rect 60 -595 85 -570
rect -60 -690 -40 -665
rect -20 -690 0 -665
rect 20 -690 40 -665
rect 60 -690 85 -665
rect -60 -785 -40 -760
rect -20 -785 0 -760
rect 20 -785 40 -760
rect 60 -785 85 -760
rect -60 -880 -40 -855
rect -20 -880 0 -855
rect 20 -880 40 -855
rect 60 -880 85 -855
rect -60 -975 -40 -950
rect -20 -975 0 -950
rect 20 -975 40 -950
rect 60 -975 85 -950
rect -60 -1070 -40 -1045
rect -20 -1070 0 -1045
rect 20 -1070 40 -1045
rect 60 -1070 85 -1045
rect -60 -1165 -40 -1140
rect -20 -1165 0 -1140
rect 20 -1165 40 -1140
rect 60 -1165 85 -1140
rect -60 -1260 -40 -1235
rect -20 -1260 0 -1235
rect 20 -1260 40 -1235
rect 60 -1260 85 -1235
rect -60 -1355 -40 -1330
rect -20 -1355 0 -1330
rect 20 -1355 40 -1330
rect 60 -1355 85 -1330
rect -60 -1450 -40 -1425
rect -20 -1450 0 -1425
rect 20 -1450 40 -1425
rect 60 -1450 85 -1425
rect -60 -1545 -40 -1520
rect -20 -1545 0 -1520
rect 20 -1545 40 -1520
rect 60 -1545 85 -1520
rect -60 -1640 -40 -1615
rect -20 -1640 0 -1615
rect 20 -1640 40 -1615
rect 60 -1640 85 -1615
rect -60 -1735 -40 -1710
rect -20 -1735 0 -1710
rect 20 -1735 40 -1710
rect 60 -1735 85 -1710
rect -60 -1830 -40 -1805
rect -20 -1830 0 -1805
rect 20 -1830 40 -1805
rect 60 -1830 85 -1805
rect -60 -1925 -40 -1900
rect -20 -1925 0 -1900
rect 20 -1925 40 -1900
rect 60 -1925 85 -1900
rect -60 -2020 -40 -1995
rect -20 -2020 0 -1995
rect 20 -2020 40 -1995
rect 60 -2020 85 -1995
rect -60 -2115 -40 -2090
rect -20 -2115 0 -2090
rect 20 -2115 40 -2090
rect 60 -2115 85 -2090
rect -60 -2210 -40 -2185
rect -20 -2210 0 -2185
rect 20 -2210 40 -2185
rect 60 -2210 85 -2185
rect -60 -2305 -40 -2280
rect -20 -2305 0 -2280
rect 20 -2305 40 -2280
rect 60 -2305 85 -2280
rect -60 -2400 -40 -2375
rect -20 -2400 0 -2375
rect 20 -2400 40 -2375
rect 60 -2400 85 -2375
rect -60 -2495 -40 -2470
rect -20 -2495 0 -2470
rect 20 -2495 40 -2470
rect 60 -2495 85 -2470
<< locali >>
rect 175 2365 2675 2375
rect 175 2345 200 2365
rect 220 2345 240 2365
rect 260 2345 280 2365
rect 300 2345 320 2365
rect 340 2345 360 2365
rect 380 2345 400 2365
rect 420 2345 440 2365
rect 460 2345 480 2365
rect 500 2345 520 2365
rect 540 2345 560 2365
rect 580 2345 600 2365
rect 620 2345 640 2365
rect 660 2345 680 2365
rect 700 2345 720 2365
rect 740 2345 760 2365
rect 780 2345 800 2365
rect 820 2345 840 2365
rect 860 2345 880 2365
rect 900 2345 920 2365
rect 940 2345 960 2365
rect 980 2345 1000 2365
rect 1020 2345 1040 2365
rect 1060 2345 1080 2365
rect 1100 2345 1120 2365
rect 1140 2345 1160 2365
rect 1180 2345 1200 2365
rect 1220 2345 1240 2365
rect 1260 2345 1280 2365
rect 1300 2345 1320 2365
rect 1340 2345 1360 2365
rect 1380 2345 1400 2365
rect 1420 2345 1440 2365
rect 1460 2345 1480 2365
rect 1500 2345 1520 2365
rect 1540 2345 1560 2365
rect 1580 2345 1600 2365
rect 1620 2345 1640 2365
rect 1660 2345 1680 2365
rect 1700 2345 1720 2365
rect 1740 2345 1760 2365
rect 1780 2345 1800 2365
rect 1820 2345 1840 2365
rect 1860 2345 1880 2365
rect 1900 2345 1920 2365
rect 1940 2345 1960 2365
rect 1980 2345 2000 2365
rect 2020 2345 2040 2365
rect 2060 2345 2080 2365
rect 2100 2345 2120 2365
rect 2140 2345 2160 2365
rect 2180 2345 2200 2365
rect 2220 2345 2240 2365
rect 2260 2345 2280 2365
rect 2300 2345 2320 2365
rect 2340 2345 2360 2365
rect 2380 2345 2400 2365
rect 2420 2345 2440 2365
rect 2460 2345 2480 2365
rect 2500 2345 2520 2365
rect 2540 2345 2560 2365
rect 2580 2345 2600 2365
rect 2620 2345 2640 2365
rect 2660 2345 2675 2365
rect 175 2335 2675 2345
rect 175 2297 2675 2307
rect 175 2277 200 2297
rect 220 2277 240 2297
rect 260 2277 280 2297
rect 300 2277 320 2297
rect 340 2277 360 2297
rect 380 2277 400 2297
rect 420 2277 440 2297
rect 460 2277 480 2297
rect 500 2277 520 2297
rect 540 2277 560 2297
rect 580 2277 600 2297
rect 620 2277 640 2297
rect 660 2277 680 2297
rect 700 2277 720 2297
rect 740 2277 760 2297
rect 780 2277 800 2297
rect 820 2277 840 2297
rect 860 2277 880 2297
rect 900 2277 920 2297
rect 940 2277 960 2297
rect 980 2277 1000 2297
rect 1020 2277 1040 2297
rect 1060 2277 1080 2297
rect 1100 2277 1120 2297
rect 1140 2277 1160 2297
rect 1180 2277 1200 2297
rect 1220 2277 1240 2297
rect 1260 2277 1280 2297
rect 1300 2277 1320 2297
rect 1340 2277 1360 2297
rect 1380 2277 1400 2297
rect 1420 2277 1440 2297
rect 1460 2277 1480 2297
rect 1500 2277 1520 2297
rect 1540 2277 1560 2297
rect 1580 2277 1600 2297
rect 1620 2277 1640 2297
rect 1660 2277 1680 2297
rect 1700 2277 1720 2297
rect 1740 2277 1760 2297
rect 1780 2277 1800 2297
rect 1820 2277 1840 2297
rect 1860 2277 1880 2297
rect 1900 2277 1920 2297
rect 1940 2277 1960 2297
rect 1980 2277 2000 2297
rect 2020 2277 2040 2297
rect 2060 2277 2080 2297
rect 2100 2277 2120 2297
rect 2140 2277 2160 2297
rect 2180 2277 2200 2297
rect 2220 2277 2240 2297
rect 2260 2277 2280 2297
rect 2300 2277 2320 2297
rect 2340 2277 2360 2297
rect 2380 2277 2400 2297
rect 2420 2277 2440 2297
rect 2460 2277 2480 2297
rect 2500 2277 2520 2297
rect 2540 2277 2560 2297
rect 2580 2277 2600 2297
rect 2620 2277 2640 2297
rect 2660 2277 2675 2297
rect 175 2267 2675 2277
rect 0 2255 155 2265
rect 0 2235 10 2255
rect 30 2235 50 2255
rect 70 2235 90 2255
rect 110 2235 130 2255
rect 0 2225 155 2235
rect 175 2215 2675 2225
rect 175 2195 200 2215
rect 220 2195 240 2215
rect 260 2195 280 2215
rect 300 2195 320 2215
rect 340 2195 360 2215
rect 380 2195 400 2215
rect 420 2195 440 2215
rect 460 2195 480 2215
rect 500 2195 520 2215
rect 540 2195 560 2215
rect 580 2195 600 2215
rect 620 2195 640 2215
rect 660 2195 680 2215
rect 700 2195 720 2215
rect 740 2195 760 2215
rect 780 2195 800 2215
rect 820 2195 840 2215
rect 860 2195 880 2215
rect 900 2195 920 2215
rect 940 2195 960 2215
rect 980 2195 1000 2215
rect 1020 2195 1040 2215
rect 1060 2195 1080 2215
rect 1100 2195 1120 2215
rect 1140 2195 1160 2215
rect 1180 2195 1200 2215
rect 1220 2195 1240 2215
rect 1260 2195 1280 2215
rect 1300 2195 1320 2215
rect 1340 2195 1360 2215
rect 1380 2195 1400 2215
rect 1420 2195 1440 2215
rect 1460 2195 1480 2215
rect 1500 2195 1520 2215
rect 1540 2195 1560 2215
rect 1580 2195 1600 2215
rect 1620 2195 1640 2215
rect 1660 2195 1680 2215
rect 1700 2195 1720 2215
rect 1740 2195 1760 2215
rect 1780 2195 1800 2215
rect 1820 2195 1840 2215
rect 1860 2195 1880 2215
rect 1900 2195 1920 2215
rect 1940 2195 1960 2215
rect 1980 2195 2000 2215
rect 2020 2195 2040 2215
rect 2060 2195 2080 2215
rect 2100 2195 2120 2215
rect 2140 2195 2160 2215
rect 2180 2195 2200 2215
rect 2220 2195 2240 2215
rect 2260 2195 2280 2215
rect 2300 2195 2320 2215
rect 2340 2195 2360 2215
rect 2380 2195 2400 2215
rect 2420 2195 2440 2215
rect 2460 2195 2480 2215
rect 2500 2195 2520 2215
rect 2540 2195 2560 2215
rect 2580 2195 2600 2215
rect 2620 2195 2640 2215
rect 2660 2195 2675 2215
rect 175 2185 2675 2195
rect 0 2175 155 2185
rect 0 2155 10 2175
rect 30 2155 50 2175
rect 70 2155 90 2175
rect 110 2155 130 2175
rect 0 2145 155 2155
rect 175 2133 2675 2143
rect 175 2113 200 2133
rect 220 2113 240 2133
rect 260 2113 280 2133
rect 300 2113 320 2133
rect 340 2113 360 2133
rect 380 2113 400 2133
rect 420 2113 440 2133
rect 460 2113 480 2133
rect 500 2113 520 2133
rect 540 2113 560 2133
rect 580 2113 600 2133
rect 620 2113 640 2133
rect 660 2113 680 2133
rect 700 2113 720 2133
rect 740 2113 760 2133
rect 780 2113 800 2133
rect 820 2113 840 2133
rect 860 2113 880 2133
rect 900 2113 920 2133
rect 940 2113 960 2133
rect 980 2113 1000 2133
rect 1020 2113 1040 2133
rect 1060 2113 1080 2133
rect 1100 2113 1120 2133
rect 1140 2113 1160 2133
rect 1180 2113 1200 2133
rect 1220 2113 1240 2133
rect 1260 2113 1280 2133
rect 1300 2113 1320 2133
rect 1340 2113 1360 2133
rect 1380 2113 1400 2133
rect 1420 2113 1440 2133
rect 1460 2113 1480 2133
rect 1500 2113 1520 2133
rect 1540 2113 1560 2133
rect 1580 2113 1600 2133
rect 1620 2113 1640 2133
rect 1660 2113 1680 2133
rect 1700 2113 1720 2133
rect 1740 2113 1760 2133
rect 1780 2113 1800 2133
rect 1820 2113 1840 2133
rect 1860 2113 1880 2133
rect 1900 2113 1920 2133
rect 1940 2113 1960 2133
rect 1980 2113 2000 2133
rect 2020 2113 2040 2133
rect 2060 2113 2080 2133
rect 2100 2113 2120 2133
rect 2140 2113 2160 2133
rect 2180 2113 2200 2133
rect 2220 2113 2240 2133
rect 2260 2113 2280 2133
rect 2300 2113 2320 2133
rect 2340 2113 2360 2133
rect 2380 2113 2400 2133
rect 2420 2113 2440 2133
rect 2460 2113 2480 2133
rect 2500 2113 2520 2133
rect 2540 2113 2560 2133
rect 2580 2113 2600 2133
rect 2620 2113 2640 2133
rect 2660 2113 2675 2133
rect 175 2103 2675 2113
rect 0 2090 155 2100
rect 0 2070 10 2090
rect 30 2070 50 2090
rect 70 2070 90 2090
rect 110 2070 130 2090
rect 0 2060 155 2070
rect 175 2051 2675 2061
rect 175 2031 200 2051
rect 220 2031 240 2051
rect 260 2031 280 2051
rect 300 2031 320 2051
rect 340 2031 360 2051
rect 380 2031 400 2051
rect 420 2031 440 2051
rect 460 2031 480 2051
rect 500 2031 520 2051
rect 540 2031 560 2051
rect 580 2031 600 2051
rect 620 2031 640 2051
rect 660 2031 680 2051
rect 700 2031 720 2051
rect 740 2031 760 2051
rect 780 2031 800 2051
rect 820 2031 840 2051
rect 860 2031 880 2051
rect 900 2031 920 2051
rect 940 2031 960 2051
rect 980 2031 1000 2051
rect 1020 2031 1040 2051
rect 1060 2031 1080 2051
rect 1100 2031 1120 2051
rect 1140 2031 1160 2051
rect 1180 2031 1200 2051
rect 1220 2031 1240 2051
rect 1260 2031 1280 2051
rect 1300 2031 1320 2051
rect 1340 2031 1360 2051
rect 1380 2031 1400 2051
rect 1420 2031 1440 2051
rect 1460 2031 1480 2051
rect 1500 2031 1520 2051
rect 1540 2031 1560 2051
rect 1580 2031 1600 2051
rect 1620 2031 1640 2051
rect 1660 2031 1680 2051
rect 1700 2031 1720 2051
rect 1740 2031 1760 2051
rect 1780 2031 1800 2051
rect 1820 2031 1840 2051
rect 1860 2031 1880 2051
rect 1900 2031 1920 2051
rect 1940 2031 1960 2051
rect 1980 2031 2000 2051
rect 2020 2031 2040 2051
rect 2060 2031 2080 2051
rect 2100 2031 2120 2051
rect 2140 2031 2160 2051
rect 2180 2031 2200 2051
rect 2220 2031 2240 2051
rect 2260 2031 2280 2051
rect 2300 2031 2320 2051
rect 2340 2031 2360 2051
rect 2380 2031 2400 2051
rect 2420 2031 2440 2051
rect 2460 2031 2480 2051
rect 2500 2031 2520 2051
rect 2540 2031 2560 2051
rect 2580 2031 2600 2051
rect 2620 2031 2640 2051
rect 2660 2031 2675 2051
rect 175 2021 2675 2031
rect 0 2010 155 2020
rect 0 1990 10 2010
rect 30 1990 50 2010
rect 70 1990 90 2010
rect 110 1990 130 2010
rect 0 1980 155 1990
rect 175 1969 2675 1979
rect 175 1949 200 1969
rect 220 1949 240 1969
rect 260 1949 280 1969
rect 300 1949 320 1969
rect 340 1949 360 1969
rect 380 1949 400 1969
rect 420 1949 440 1969
rect 460 1949 480 1969
rect 500 1949 520 1969
rect 540 1949 560 1969
rect 580 1949 600 1969
rect 620 1949 640 1969
rect 660 1949 680 1969
rect 700 1949 720 1969
rect 740 1949 760 1969
rect 780 1949 800 1969
rect 820 1949 840 1969
rect 860 1949 880 1969
rect 900 1949 920 1969
rect 940 1949 960 1969
rect 980 1949 1000 1969
rect 1020 1949 1040 1969
rect 1060 1949 1080 1969
rect 1100 1949 1120 1969
rect 1140 1949 1160 1969
rect 1180 1949 1200 1969
rect 1220 1949 1240 1969
rect 1260 1949 1280 1969
rect 1300 1949 1320 1969
rect 1340 1949 1360 1969
rect 1380 1949 1400 1969
rect 1420 1949 1440 1969
rect 1460 1949 1480 1969
rect 1500 1949 1520 1969
rect 1540 1949 1560 1969
rect 1580 1949 1600 1969
rect 1620 1949 1640 1969
rect 1660 1949 1680 1969
rect 1700 1949 1720 1969
rect 1740 1949 1760 1969
rect 1780 1949 1800 1969
rect 1820 1949 1840 1969
rect 1860 1949 1880 1969
rect 1900 1949 1920 1969
rect 1940 1949 1960 1969
rect 1980 1949 2000 1969
rect 2020 1949 2040 1969
rect 2060 1949 2080 1969
rect 2100 1949 2120 1969
rect 2140 1949 2160 1969
rect 2180 1949 2200 1969
rect 2220 1949 2240 1969
rect 2260 1949 2280 1969
rect 2300 1949 2320 1969
rect 2340 1949 2360 1969
rect 2380 1949 2400 1969
rect 2420 1949 2440 1969
rect 2460 1949 2480 1969
rect 2500 1949 2520 1969
rect 2540 1949 2560 1969
rect 2580 1949 2600 1969
rect 2620 1949 2640 1969
rect 2660 1949 2675 1969
rect 0 1930 155 1940
rect 175 1939 2675 1949
rect 0 1910 10 1930
rect 30 1910 50 1930
rect 70 1910 90 1930
rect 110 1910 130 1930
rect 0 1900 155 1910
rect 175 1887 2675 1897
rect 175 1867 200 1887
rect 220 1867 240 1887
rect 260 1867 280 1887
rect 300 1867 320 1887
rect 340 1867 360 1887
rect 380 1867 400 1887
rect 420 1867 440 1887
rect 460 1867 480 1887
rect 500 1867 520 1887
rect 540 1867 560 1887
rect 580 1867 600 1887
rect 620 1867 640 1887
rect 660 1867 680 1887
rect 700 1867 720 1887
rect 740 1867 760 1887
rect 780 1867 800 1887
rect 820 1867 840 1887
rect 860 1867 880 1887
rect 900 1867 920 1887
rect 940 1867 960 1887
rect 980 1867 1000 1887
rect 1020 1867 1040 1887
rect 1060 1867 1080 1887
rect 1100 1867 1120 1887
rect 1140 1867 1160 1887
rect 1180 1867 1200 1887
rect 1220 1867 1240 1887
rect 1260 1867 1280 1887
rect 1300 1867 1320 1887
rect 1340 1867 1360 1887
rect 1380 1867 1400 1887
rect 1420 1867 1440 1887
rect 1460 1867 1480 1887
rect 1500 1867 1520 1887
rect 1540 1867 1560 1887
rect 1580 1867 1600 1887
rect 1620 1867 1640 1887
rect 1660 1867 1680 1887
rect 1700 1867 1720 1887
rect 1740 1867 1760 1887
rect 1780 1867 1800 1887
rect 1820 1867 1840 1887
rect 1860 1867 1880 1887
rect 1900 1867 1920 1887
rect 1940 1867 1960 1887
rect 1980 1867 2000 1887
rect 2020 1867 2040 1887
rect 2060 1867 2080 1887
rect 2100 1867 2120 1887
rect 2140 1867 2160 1887
rect 2180 1867 2200 1887
rect 2220 1867 2240 1887
rect 2260 1867 2280 1887
rect 2300 1867 2320 1887
rect 2340 1867 2360 1887
rect 2380 1867 2400 1887
rect 2420 1867 2440 1887
rect 2460 1867 2480 1887
rect 2500 1867 2520 1887
rect 2540 1867 2560 1887
rect 2580 1867 2600 1887
rect 2620 1867 2640 1887
rect 2660 1867 2675 1887
rect 175 1857 2675 1867
rect 0 1845 155 1855
rect 0 1825 10 1845
rect 30 1825 50 1845
rect 70 1825 90 1845
rect 110 1825 130 1845
rect 0 1815 155 1825
rect 175 1805 2675 1815
rect 175 1785 200 1805
rect 220 1785 240 1805
rect 260 1785 280 1805
rect 300 1785 320 1805
rect 340 1785 360 1805
rect 380 1785 400 1805
rect 420 1785 440 1805
rect 460 1785 480 1805
rect 500 1785 520 1805
rect 540 1785 560 1805
rect 580 1785 600 1805
rect 620 1785 640 1805
rect 660 1785 680 1805
rect 700 1785 720 1805
rect 740 1785 760 1805
rect 780 1785 800 1805
rect 820 1785 840 1805
rect 860 1785 880 1805
rect 900 1785 920 1805
rect 940 1785 960 1805
rect 980 1785 1000 1805
rect 1020 1785 1040 1805
rect 1060 1785 1080 1805
rect 1100 1785 1120 1805
rect 1140 1785 1160 1805
rect 1180 1785 1200 1805
rect 1220 1785 1240 1805
rect 1260 1785 1280 1805
rect 1300 1785 1320 1805
rect 1340 1785 1360 1805
rect 1380 1785 1400 1805
rect 1420 1785 1440 1805
rect 1460 1785 1480 1805
rect 1500 1785 1520 1805
rect 1540 1785 1560 1805
rect 1580 1785 1600 1805
rect 1620 1785 1640 1805
rect 1660 1785 1680 1805
rect 1700 1785 1720 1805
rect 1740 1785 1760 1805
rect 1780 1785 1800 1805
rect 1820 1785 1840 1805
rect 1860 1785 1880 1805
rect 1900 1785 1920 1805
rect 1940 1785 1960 1805
rect 1980 1785 2000 1805
rect 2020 1785 2040 1805
rect 2060 1785 2080 1805
rect 2100 1785 2120 1805
rect 2140 1785 2160 1805
rect 2180 1785 2200 1805
rect 2220 1785 2240 1805
rect 2260 1785 2280 1805
rect 2300 1785 2320 1805
rect 2340 1785 2360 1805
rect 2380 1785 2400 1805
rect 2420 1785 2440 1805
rect 2460 1785 2480 1805
rect 2500 1785 2520 1805
rect 2540 1785 2560 1805
rect 2580 1785 2600 1805
rect 2620 1785 2640 1805
rect 2660 1785 2675 1805
rect 175 1775 2675 1785
rect 0 1765 155 1775
rect 0 1745 10 1765
rect 30 1745 50 1765
rect 70 1745 90 1765
rect 110 1745 130 1765
rect 0 1735 155 1745
rect 175 1723 2675 1733
rect 175 1703 200 1723
rect 220 1703 240 1723
rect 260 1703 280 1723
rect 300 1703 320 1723
rect 340 1703 360 1723
rect 380 1703 400 1723
rect 420 1703 440 1723
rect 460 1703 480 1723
rect 500 1703 520 1723
rect 540 1703 560 1723
rect 580 1703 600 1723
rect 620 1703 640 1723
rect 660 1703 680 1723
rect 700 1703 720 1723
rect 740 1703 760 1723
rect 780 1703 800 1723
rect 820 1703 840 1723
rect 860 1703 880 1723
rect 900 1703 920 1723
rect 940 1703 960 1723
rect 980 1703 1000 1723
rect 1020 1703 1040 1723
rect 1060 1703 1080 1723
rect 1100 1703 1120 1723
rect 1140 1703 1160 1723
rect 1180 1703 1200 1723
rect 1220 1703 1240 1723
rect 1260 1703 1280 1723
rect 1300 1703 1320 1723
rect 1340 1703 1360 1723
rect 1380 1703 1400 1723
rect 1420 1703 1440 1723
rect 1460 1703 1480 1723
rect 1500 1703 1520 1723
rect 1540 1703 1560 1723
rect 1580 1703 1600 1723
rect 1620 1703 1640 1723
rect 1660 1703 1680 1723
rect 1700 1703 1720 1723
rect 1740 1703 1760 1723
rect 1780 1703 1800 1723
rect 1820 1703 1840 1723
rect 1860 1703 1880 1723
rect 1900 1703 1920 1723
rect 1940 1703 1960 1723
rect 1980 1703 2000 1723
rect 2020 1703 2040 1723
rect 2060 1703 2080 1723
rect 2100 1703 2120 1723
rect 2140 1703 2160 1723
rect 2180 1703 2200 1723
rect 2220 1703 2240 1723
rect 2260 1703 2280 1723
rect 2300 1703 2320 1723
rect 2340 1703 2360 1723
rect 2380 1703 2400 1723
rect 2420 1703 2440 1723
rect 2460 1703 2480 1723
rect 2500 1703 2520 1723
rect 2540 1703 2560 1723
rect 2580 1703 2600 1723
rect 2620 1703 2640 1723
rect 2660 1703 2675 1723
rect 175 1693 2675 1703
rect 0 1680 155 1690
rect 0 1660 10 1680
rect 30 1660 50 1680
rect 70 1660 90 1680
rect 110 1660 130 1680
rect 0 1650 155 1660
rect 175 1641 2675 1651
rect 175 1621 200 1641
rect 220 1621 240 1641
rect 260 1621 280 1641
rect 300 1621 320 1641
rect 340 1621 360 1641
rect 380 1621 400 1641
rect 420 1621 440 1641
rect 460 1621 480 1641
rect 500 1621 520 1641
rect 540 1621 560 1641
rect 580 1621 600 1641
rect 620 1621 640 1641
rect 660 1621 680 1641
rect 700 1621 720 1641
rect 740 1621 760 1641
rect 780 1621 800 1641
rect 820 1621 840 1641
rect 860 1621 880 1641
rect 900 1621 920 1641
rect 940 1621 960 1641
rect 980 1621 1000 1641
rect 1020 1621 1040 1641
rect 1060 1621 1080 1641
rect 1100 1621 1120 1641
rect 1140 1621 1160 1641
rect 1180 1621 1200 1641
rect 1220 1621 1240 1641
rect 1260 1621 1280 1641
rect 1300 1621 1320 1641
rect 1340 1621 1360 1641
rect 1380 1621 1400 1641
rect 1420 1621 1440 1641
rect 1460 1621 1480 1641
rect 1500 1621 1520 1641
rect 1540 1621 1560 1641
rect 1580 1621 1600 1641
rect 1620 1621 1640 1641
rect 1660 1621 1680 1641
rect 1700 1621 1720 1641
rect 1740 1621 1760 1641
rect 1780 1621 1800 1641
rect 1820 1621 1840 1641
rect 1860 1621 1880 1641
rect 1900 1621 1920 1641
rect 1940 1621 1960 1641
rect 1980 1621 2000 1641
rect 2020 1621 2040 1641
rect 2060 1621 2080 1641
rect 2100 1621 2120 1641
rect 2140 1621 2160 1641
rect 2180 1621 2200 1641
rect 2220 1621 2240 1641
rect 2260 1621 2280 1641
rect 2300 1621 2320 1641
rect 2340 1621 2360 1641
rect 2380 1621 2400 1641
rect 2420 1621 2440 1641
rect 2460 1621 2480 1641
rect 2500 1621 2520 1641
rect 2540 1621 2560 1641
rect 2580 1621 2600 1641
rect 2620 1621 2640 1641
rect 2660 1621 2675 1641
rect 175 1611 2675 1621
rect 0 1600 155 1610
rect 0 1580 10 1600
rect 30 1580 50 1600
rect 70 1580 90 1600
rect 110 1580 130 1600
rect 0 1570 155 1580
rect 175 1559 2675 1569
rect 175 1539 200 1559
rect 220 1539 240 1559
rect 260 1539 280 1559
rect 300 1539 320 1559
rect 340 1539 360 1559
rect 380 1539 400 1559
rect 420 1539 440 1559
rect 460 1539 480 1559
rect 500 1539 520 1559
rect 540 1539 560 1559
rect 580 1539 600 1559
rect 620 1539 640 1559
rect 660 1539 680 1559
rect 700 1539 720 1559
rect 740 1539 760 1559
rect 780 1539 800 1559
rect 820 1539 840 1559
rect 860 1539 880 1559
rect 900 1539 920 1559
rect 940 1539 960 1559
rect 980 1539 1000 1559
rect 1020 1539 1040 1559
rect 1060 1539 1080 1559
rect 1100 1539 1120 1559
rect 1140 1539 1160 1559
rect 1180 1539 1200 1559
rect 1220 1539 1240 1559
rect 1260 1539 1280 1559
rect 1300 1539 1320 1559
rect 1340 1539 1360 1559
rect 1380 1539 1400 1559
rect 1420 1539 1440 1559
rect 1460 1539 1480 1559
rect 1500 1539 1520 1559
rect 1540 1539 1560 1559
rect 1580 1539 1600 1559
rect 1620 1539 1640 1559
rect 1660 1539 1680 1559
rect 1700 1539 1720 1559
rect 1740 1539 1760 1559
rect 1780 1539 1800 1559
rect 1820 1539 1840 1559
rect 1860 1539 1880 1559
rect 1900 1539 1920 1559
rect 1940 1539 1960 1559
rect 1980 1539 2000 1559
rect 2020 1539 2040 1559
rect 2060 1539 2080 1559
rect 2100 1539 2120 1559
rect 2140 1539 2160 1559
rect 2180 1539 2200 1559
rect 2220 1539 2240 1559
rect 2260 1539 2280 1559
rect 2300 1539 2320 1559
rect 2340 1539 2360 1559
rect 2380 1539 2400 1559
rect 2420 1539 2440 1559
rect 2460 1539 2480 1559
rect 2500 1539 2520 1559
rect 2540 1539 2560 1559
rect 2580 1539 2600 1559
rect 2620 1539 2640 1559
rect 2660 1539 2675 1559
rect 0 1520 155 1530
rect 175 1529 2675 1539
rect 0 1500 10 1520
rect 30 1500 50 1520
rect 70 1500 90 1520
rect 110 1500 130 1520
rect 0 1490 155 1500
rect 175 1477 2675 1487
rect 175 1457 200 1477
rect 220 1457 240 1477
rect 260 1457 280 1477
rect 300 1457 320 1477
rect 340 1457 360 1477
rect 380 1457 400 1477
rect 420 1457 440 1477
rect 460 1457 480 1477
rect 500 1457 520 1477
rect 540 1457 560 1477
rect 580 1457 600 1477
rect 620 1457 640 1477
rect 660 1457 680 1477
rect 700 1457 720 1477
rect 740 1457 760 1477
rect 780 1457 800 1477
rect 820 1457 840 1477
rect 860 1457 880 1477
rect 900 1457 920 1477
rect 940 1457 960 1477
rect 980 1457 1000 1477
rect 1020 1457 1040 1477
rect 1060 1457 1080 1477
rect 1100 1457 1120 1477
rect 1140 1457 1160 1477
rect 1180 1457 1200 1477
rect 1220 1457 1240 1477
rect 1260 1457 1280 1477
rect 1300 1457 1320 1477
rect 1340 1457 1360 1477
rect 1380 1457 1400 1477
rect 1420 1457 1440 1477
rect 1460 1457 1480 1477
rect 1500 1457 1520 1477
rect 1540 1457 1560 1477
rect 1580 1457 1600 1477
rect 1620 1457 1640 1477
rect 1660 1457 1680 1477
rect 1700 1457 1720 1477
rect 1740 1457 1760 1477
rect 1780 1457 1800 1477
rect 1820 1457 1840 1477
rect 1860 1457 1880 1477
rect 1900 1457 1920 1477
rect 1940 1457 1960 1477
rect 1980 1457 2000 1477
rect 2020 1457 2040 1477
rect 2060 1457 2080 1477
rect 2100 1457 2120 1477
rect 2140 1457 2160 1477
rect 2180 1457 2200 1477
rect 2220 1457 2240 1477
rect 2260 1457 2280 1477
rect 2300 1457 2320 1477
rect 2340 1457 2360 1477
rect 2380 1457 2400 1477
rect 2420 1457 2440 1477
rect 2460 1457 2480 1477
rect 2500 1457 2520 1477
rect 2540 1457 2560 1477
rect 2580 1457 2600 1477
rect 2620 1457 2640 1477
rect 2660 1457 2675 1477
rect 175 1447 2675 1457
rect 0 1435 155 1445
rect 0 1415 10 1435
rect 30 1415 50 1435
rect 70 1415 90 1435
rect 110 1415 130 1435
rect 0 1405 155 1415
rect 175 1395 2675 1405
rect 175 1375 200 1395
rect 220 1375 240 1395
rect 260 1375 280 1395
rect 300 1375 320 1395
rect 340 1375 360 1395
rect 380 1375 400 1395
rect 420 1375 440 1395
rect 460 1375 480 1395
rect 500 1375 520 1395
rect 540 1375 560 1395
rect 580 1375 600 1395
rect 620 1375 640 1395
rect 660 1375 680 1395
rect 700 1375 720 1395
rect 740 1375 760 1395
rect 780 1375 800 1395
rect 820 1375 840 1395
rect 860 1375 880 1395
rect 900 1375 920 1395
rect 940 1375 960 1395
rect 980 1375 1000 1395
rect 1020 1375 1040 1395
rect 1060 1375 1080 1395
rect 1100 1375 1120 1395
rect 1140 1375 1160 1395
rect 1180 1375 1200 1395
rect 1220 1375 1240 1395
rect 1260 1375 1280 1395
rect 1300 1375 1320 1395
rect 1340 1375 1360 1395
rect 1380 1375 1400 1395
rect 1420 1375 1440 1395
rect 1460 1375 1480 1395
rect 1500 1375 1520 1395
rect 1540 1375 1560 1395
rect 1580 1375 1600 1395
rect 1620 1375 1640 1395
rect 1660 1375 1680 1395
rect 1700 1375 1720 1395
rect 1740 1375 1760 1395
rect 1780 1375 1800 1395
rect 1820 1375 1840 1395
rect 1860 1375 1880 1395
rect 1900 1375 1920 1395
rect 1940 1375 1960 1395
rect 1980 1375 2000 1395
rect 2020 1375 2040 1395
rect 2060 1375 2080 1395
rect 2100 1375 2120 1395
rect 2140 1375 2160 1395
rect 2180 1375 2200 1395
rect 2220 1375 2240 1395
rect 2260 1375 2280 1395
rect 2300 1375 2320 1395
rect 2340 1375 2360 1395
rect 2380 1375 2400 1395
rect 2420 1375 2440 1395
rect 2460 1375 2480 1395
rect 2500 1375 2520 1395
rect 2540 1375 2560 1395
rect 2580 1375 2600 1395
rect 2620 1375 2640 1395
rect 2660 1375 2675 1395
rect 175 1365 2675 1375
rect 0 1355 155 1365
rect 0 1335 10 1355
rect 30 1335 50 1355
rect 70 1335 90 1355
rect 110 1335 130 1355
rect 0 1325 155 1335
rect 175 1313 2675 1323
rect 175 1293 200 1313
rect 220 1293 240 1313
rect 260 1293 280 1313
rect 300 1293 320 1313
rect 340 1293 360 1313
rect 380 1293 400 1313
rect 420 1293 440 1313
rect 460 1293 480 1313
rect 500 1293 520 1313
rect 540 1293 560 1313
rect 580 1293 600 1313
rect 620 1293 640 1313
rect 660 1293 680 1313
rect 700 1293 720 1313
rect 740 1293 760 1313
rect 780 1293 800 1313
rect 820 1293 840 1313
rect 860 1293 880 1313
rect 900 1293 920 1313
rect 940 1293 960 1313
rect 980 1293 1000 1313
rect 1020 1293 1040 1313
rect 1060 1293 1080 1313
rect 1100 1293 1120 1313
rect 1140 1293 1160 1313
rect 1180 1293 1200 1313
rect 1220 1293 1240 1313
rect 1260 1293 1280 1313
rect 1300 1293 1320 1313
rect 1340 1293 1360 1313
rect 1380 1293 1400 1313
rect 1420 1293 1440 1313
rect 1460 1293 1480 1313
rect 1500 1293 1520 1313
rect 1540 1293 1560 1313
rect 1580 1293 1600 1313
rect 1620 1293 1640 1313
rect 1660 1293 1680 1313
rect 1700 1293 1720 1313
rect 1740 1293 1760 1313
rect 1780 1293 1800 1313
rect 1820 1293 1840 1313
rect 1860 1293 1880 1313
rect 1900 1293 1920 1313
rect 1940 1293 1960 1313
rect 1980 1293 2000 1313
rect 2020 1293 2040 1313
rect 2060 1293 2080 1313
rect 2100 1293 2120 1313
rect 2140 1293 2160 1313
rect 2180 1293 2200 1313
rect 2220 1293 2240 1313
rect 2260 1293 2280 1313
rect 2300 1293 2320 1313
rect 2340 1293 2360 1313
rect 2380 1293 2400 1313
rect 2420 1293 2440 1313
rect 2460 1293 2480 1313
rect 2500 1293 2520 1313
rect 2540 1293 2560 1313
rect 2580 1293 2600 1313
rect 2620 1293 2640 1313
rect 2660 1293 2675 1313
rect 175 1283 2675 1293
rect 0 1270 155 1280
rect 0 1250 10 1270
rect 30 1250 50 1270
rect 70 1250 90 1270
rect 110 1250 130 1270
rect 0 1240 155 1250
rect 175 1231 2675 1241
rect 175 1211 200 1231
rect 220 1211 240 1231
rect 260 1211 280 1231
rect 300 1211 320 1231
rect 340 1211 360 1231
rect 380 1211 400 1231
rect 420 1211 440 1231
rect 460 1211 480 1231
rect 500 1211 520 1231
rect 540 1211 560 1231
rect 580 1211 600 1231
rect 620 1211 640 1231
rect 660 1211 680 1231
rect 700 1211 720 1231
rect 740 1211 760 1231
rect 780 1211 800 1231
rect 820 1211 840 1231
rect 860 1211 880 1231
rect 900 1211 920 1231
rect 940 1211 960 1231
rect 980 1211 1000 1231
rect 1020 1211 1040 1231
rect 1060 1211 1080 1231
rect 1100 1211 1120 1231
rect 1140 1211 1160 1231
rect 1180 1211 1200 1231
rect 1220 1211 1240 1231
rect 1260 1211 1280 1231
rect 1300 1211 1320 1231
rect 1340 1211 1360 1231
rect 1380 1211 1400 1231
rect 1420 1211 1440 1231
rect 1460 1211 1480 1231
rect 1500 1211 1520 1231
rect 1540 1211 1560 1231
rect 1580 1211 1600 1231
rect 1620 1211 1640 1231
rect 1660 1211 1680 1231
rect 1700 1211 1720 1231
rect 1740 1211 1760 1231
rect 1780 1211 1800 1231
rect 1820 1211 1840 1231
rect 1860 1211 1880 1231
rect 1900 1211 1920 1231
rect 1940 1211 1960 1231
rect 1980 1211 2000 1231
rect 2020 1211 2040 1231
rect 2060 1211 2080 1231
rect 2100 1211 2120 1231
rect 2140 1211 2160 1231
rect 2180 1211 2200 1231
rect 2220 1211 2240 1231
rect 2260 1211 2280 1231
rect 2300 1211 2320 1231
rect 2340 1211 2360 1231
rect 2380 1211 2400 1231
rect 2420 1211 2440 1231
rect 2460 1211 2480 1231
rect 2500 1211 2520 1231
rect 2540 1211 2560 1231
rect 2580 1211 2600 1231
rect 2620 1211 2640 1231
rect 2660 1211 2675 1231
rect 175 1201 2675 1211
rect 0 1190 155 1200
rect 0 1170 10 1190
rect 30 1170 50 1190
rect 70 1170 90 1190
rect 110 1170 130 1190
rect 0 1160 155 1170
rect 175 1149 2675 1159
rect 175 1129 200 1149
rect 220 1129 240 1149
rect 260 1129 280 1149
rect 300 1129 320 1149
rect 340 1129 360 1149
rect 380 1129 400 1149
rect 420 1129 440 1149
rect 460 1129 480 1149
rect 500 1129 520 1149
rect 540 1129 560 1149
rect 580 1129 600 1149
rect 620 1129 640 1149
rect 660 1129 680 1149
rect 700 1129 720 1149
rect 740 1129 760 1149
rect 780 1129 800 1149
rect 820 1129 840 1149
rect 860 1129 880 1149
rect 900 1129 920 1149
rect 940 1129 960 1149
rect 980 1129 1000 1149
rect 1020 1129 1040 1149
rect 1060 1129 1080 1149
rect 1100 1129 1120 1149
rect 1140 1129 1160 1149
rect 1180 1129 1200 1149
rect 1220 1129 1240 1149
rect 1260 1129 1280 1149
rect 1300 1129 1320 1149
rect 1340 1129 1360 1149
rect 1380 1129 1400 1149
rect 1420 1129 1440 1149
rect 1460 1129 1480 1149
rect 1500 1129 1520 1149
rect 1540 1129 1560 1149
rect 1580 1129 1600 1149
rect 1620 1129 1640 1149
rect 1660 1129 1680 1149
rect 1700 1129 1720 1149
rect 1740 1129 1760 1149
rect 1780 1129 1800 1149
rect 1820 1129 1840 1149
rect 1860 1129 1880 1149
rect 1900 1129 1920 1149
rect 1940 1129 1960 1149
rect 1980 1129 2000 1149
rect 2020 1129 2040 1149
rect 2060 1129 2080 1149
rect 2100 1129 2120 1149
rect 2140 1129 2160 1149
rect 2180 1129 2200 1149
rect 2220 1129 2240 1149
rect 2260 1129 2280 1149
rect 2300 1129 2320 1149
rect 2340 1129 2360 1149
rect 2380 1129 2400 1149
rect 2420 1129 2440 1149
rect 2460 1129 2480 1149
rect 2500 1129 2520 1149
rect 2540 1129 2560 1149
rect 2580 1129 2600 1149
rect 2620 1129 2640 1149
rect 2660 1129 2675 1149
rect 0 1110 155 1120
rect 175 1119 2675 1129
rect 0 1090 10 1110
rect 30 1090 50 1110
rect 70 1090 90 1110
rect 110 1090 130 1110
rect 0 1080 155 1090
rect 175 1067 2675 1077
rect 175 1047 200 1067
rect 220 1047 240 1067
rect 260 1047 280 1067
rect 300 1047 320 1067
rect 340 1047 360 1067
rect 380 1047 400 1067
rect 420 1047 440 1067
rect 460 1047 480 1067
rect 500 1047 520 1067
rect 540 1047 560 1067
rect 580 1047 600 1067
rect 620 1047 640 1067
rect 660 1047 680 1067
rect 700 1047 720 1067
rect 740 1047 760 1067
rect 780 1047 800 1067
rect 820 1047 840 1067
rect 860 1047 880 1067
rect 900 1047 920 1067
rect 940 1047 960 1067
rect 980 1047 1000 1067
rect 1020 1047 1040 1067
rect 1060 1047 1080 1067
rect 1100 1047 1120 1067
rect 1140 1047 1160 1067
rect 1180 1047 1200 1067
rect 1220 1047 1240 1067
rect 1260 1047 1280 1067
rect 1300 1047 1320 1067
rect 1340 1047 1360 1067
rect 1380 1047 1400 1067
rect 1420 1047 1440 1067
rect 1460 1047 1480 1067
rect 1500 1047 1520 1067
rect 1540 1047 1560 1067
rect 1580 1047 1600 1067
rect 1620 1047 1640 1067
rect 1660 1047 1680 1067
rect 1700 1047 1720 1067
rect 1740 1047 1760 1067
rect 1780 1047 1800 1067
rect 1820 1047 1840 1067
rect 1860 1047 1880 1067
rect 1900 1047 1920 1067
rect 1940 1047 1960 1067
rect 1980 1047 2000 1067
rect 2020 1047 2040 1067
rect 2060 1047 2080 1067
rect 2100 1047 2120 1067
rect 2140 1047 2160 1067
rect 2180 1047 2200 1067
rect 2220 1047 2240 1067
rect 2260 1047 2280 1067
rect 2300 1047 2320 1067
rect 2340 1047 2360 1067
rect 2380 1047 2400 1067
rect 2420 1047 2440 1067
rect 2460 1047 2480 1067
rect 2500 1047 2520 1067
rect 2540 1047 2560 1067
rect 2580 1047 2600 1067
rect 2620 1047 2640 1067
rect 2660 1047 2675 1067
rect 175 1037 2675 1047
rect 0 1025 155 1035
rect 0 1005 10 1025
rect 30 1005 50 1025
rect 70 1005 90 1025
rect 110 1005 130 1025
rect 0 995 155 1005
rect 175 985 2675 995
rect 175 965 200 985
rect 220 965 240 985
rect 260 965 280 985
rect 300 965 320 985
rect 340 965 360 985
rect 380 965 400 985
rect 420 965 440 985
rect 460 965 480 985
rect 500 965 520 985
rect 540 965 560 985
rect 580 965 600 985
rect 620 965 640 985
rect 660 965 680 985
rect 700 965 720 985
rect 740 965 760 985
rect 780 965 800 985
rect 820 965 840 985
rect 860 965 880 985
rect 900 965 920 985
rect 940 965 960 985
rect 980 965 1000 985
rect 1020 965 1040 985
rect 1060 965 1080 985
rect 1100 965 1120 985
rect 1140 965 1160 985
rect 1180 965 1200 985
rect 1220 965 1240 985
rect 1260 965 1280 985
rect 1300 965 1320 985
rect 1340 965 1360 985
rect 1380 965 1400 985
rect 1420 965 1440 985
rect 1460 965 1480 985
rect 1500 965 1520 985
rect 1540 965 1560 985
rect 1580 965 1600 985
rect 1620 965 1640 985
rect 1660 965 1680 985
rect 1700 965 1720 985
rect 1740 965 1760 985
rect 1780 965 1800 985
rect 1820 965 1840 985
rect 1860 965 1880 985
rect 1900 965 1920 985
rect 1940 965 1960 985
rect 1980 965 2000 985
rect 2020 965 2040 985
rect 2060 965 2080 985
rect 2100 965 2120 985
rect 2140 965 2160 985
rect 2180 965 2200 985
rect 2220 965 2240 985
rect 2260 965 2280 985
rect 2300 965 2320 985
rect 2340 965 2360 985
rect 2380 965 2400 985
rect 2420 965 2440 985
rect 2460 965 2480 985
rect 2500 965 2520 985
rect 2540 965 2560 985
rect 2580 965 2600 985
rect 2620 965 2640 985
rect 2660 965 2675 985
rect 175 955 2675 965
rect 0 945 155 955
rect 0 925 10 945
rect 30 925 50 945
rect 70 925 90 945
rect 110 925 130 945
rect 0 915 155 925
rect 175 903 2675 913
rect 175 883 200 903
rect 220 883 240 903
rect 260 883 280 903
rect 300 883 320 903
rect 340 883 360 903
rect 380 883 400 903
rect 420 883 440 903
rect 460 883 480 903
rect 500 883 520 903
rect 540 883 560 903
rect 580 883 600 903
rect 620 883 640 903
rect 660 883 680 903
rect 700 883 720 903
rect 740 883 760 903
rect 780 883 800 903
rect 820 883 840 903
rect 860 883 880 903
rect 900 883 920 903
rect 940 883 960 903
rect 980 883 1000 903
rect 1020 883 1040 903
rect 1060 883 1080 903
rect 1100 883 1120 903
rect 1140 883 1160 903
rect 1180 883 1200 903
rect 1220 883 1240 903
rect 1260 883 1280 903
rect 1300 883 1320 903
rect 1340 883 1360 903
rect 1380 883 1400 903
rect 1420 883 1440 903
rect 1460 883 1480 903
rect 1500 883 1520 903
rect 1540 883 1560 903
rect 1580 883 1600 903
rect 1620 883 1640 903
rect 1660 883 1680 903
rect 1700 883 1720 903
rect 1740 883 1760 903
rect 1780 883 1800 903
rect 1820 883 1840 903
rect 1860 883 1880 903
rect 1900 883 1920 903
rect 1940 883 1960 903
rect 1980 883 2000 903
rect 2020 883 2040 903
rect 2060 883 2080 903
rect 2100 883 2120 903
rect 2140 883 2160 903
rect 2180 883 2200 903
rect 2220 883 2240 903
rect 2260 883 2280 903
rect 2300 883 2320 903
rect 2340 883 2360 903
rect 2380 883 2400 903
rect 2420 883 2440 903
rect 2460 883 2480 903
rect 2500 883 2520 903
rect 2540 883 2560 903
rect 2580 883 2600 903
rect 2620 883 2640 903
rect 2660 883 2675 903
rect 175 873 2675 883
rect 0 860 155 870
rect 0 840 10 860
rect 30 840 50 860
rect 70 840 90 860
rect 110 840 130 860
rect 0 830 155 840
rect 175 821 2675 831
rect 175 801 200 821
rect 220 801 240 821
rect 260 801 280 821
rect 300 801 320 821
rect 340 801 360 821
rect 380 801 400 821
rect 420 801 440 821
rect 460 801 480 821
rect 500 801 520 821
rect 540 801 560 821
rect 580 801 600 821
rect 620 801 640 821
rect 660 801 680 821
rect 700 801 720 821
rect 740 801 760 821
rect 780 801 800 821
rect 820 801 840 821
rect 860 801 880 821
rect 900 801 920 821
rect 940 801 960 821
rect 980 801 1000 821
rect 1020 801 1040 821
rect 1060 801 1080 821
rect 1100 801 1120 821
rect 1140 801 1160 821
rect 1180 801 1200 821
rect 1220 801 1240 821
rect 1260 801 1280 821
rect 1300 801 1320 821
rect 1340 801 1360 821
rect 1380 801 1400 821
rect 1420 801 1440 821
rect 1460 801 1480 821
rect 1500 801 1520 821
rect 1540 801 1560 821
rect 1580 801 1600 821
rect 1620 801 1640 821
rect 1660 801 1680 821
rect 1700 801 1720 821
rect 1740 801 1760 821
rect 1780 801 1800 821
rect 1820 801 1840 821
rect 1860 801 1880 821
rect 1900 801 1920 821
rect 1940 801 1960 821
rect 1980 801 2000 821
rect 2020 801 2040 821
rect 2060 801 2080 821
rect 2100 801 2120 821
rect 2140 801 2160 821
rect 2180 801 2200 821
rect 2220 801 2240 821
rect 2260 801 2280 821
rect 2300 801 2320 821
rect 2340 801 2360 821
rect 2380 801 2400 821
rect 2420 801 2440 821
rect 2460 801 2480 821
rect 2500 801 2520 821
rect 2540 801 2560 821
rect 2580 801 2600 821
rect 2620 801 2640 821
rect 2660 801 2675 821
rect 175 791 2675 801
rect 0 780 155 790
rect 0 760 10 780
rect 30 760 50 780
rect 70 760 90 780
rect 110 760 130 780
rect 0 750 155 760
rect 175 739 2675 749
rect 175 719 200 739
rect 220 719 240 739
rect 260 719 280 739
rect 300 719 320 739
rect 340 719 360 739
rect 380 719 400 739
rect 420 719 440 739
rect 460 719 480 739
rect 500 719 520 739
rect 540 719 560 739
rect 580 719 600 739
rect 620 719 640 739
rect 660 719 680 739
rect 700 719 720 739
rect 740 719 760 739
rect 780 719 800 739
rect 820 719 840 739
rect 860 719 880 739
rect 900 719 920 739
rect 940 719 960 739
rect 980 719 1000 739
rect 1020 719 1040 739
rect 1060 719 1080 739
rect 1100 719 1120 739
rect 1140 719 1160 739
rect 1180 719 1200 739
rect 1220 719 1240 739
rect 1260 719 1280 739
rect 1300 719 1320 739
rect 1340 719 1360 739
rect 1380 719 1400 739
rect 1420 719 1440 739
rect 1460 719 1480 739
rect 1500 719 1520 739
rect 1540 719 1560 739
rect 1580 719 1600 739
rect 1620 719 1640 739
rect 1660 719 1680 739
rect 1700 719 1720 739
rect 1740 719 1760 739
rect 1780 719 1800 739
rect 1820 719 1840 739
rect 1860 719 1880 739
rect 1900 719 1920 739
rect 1940 719 1960 739
rect 1980 719 2000 739
rect 2020 719 2040 739
rect 2060 719 2080 739
rect 2100 719 2120 739
rect 2140 719 2160 739
rect 2180 719 2200 739
rect 2220 719 2240 739
rect 2260 719 2280 739
rect 2300 719 2320 739
rect 2340 719 2360 739
rect 2380 719 2400 739
rect 2420 719 2440 739
rect 2460 719 2480 739
rect 2500 719 2520 739
rect 2540 719 2560 739
rect 2580 719 2600 739
rect 2620 719 2640 739
rect 2660 719 2675 739
rect 0 700 155 710
rect 175 709 2675 719
rect 0 680 10 700
rect 30 680 50 700
rect 70 680 90 700
rect 110 680 130 700
rect 0 670 155 680
rect 175 657 2675 667
rect 175 637 200 657
rect 220 637 240 657
rect 260 637 280 657
rect 300 637 320 657
rect 340 637 360 657
rect 380 637 400 657
rect 420 637 440 657
rect 460 637 480 657
rect 500 637 520 657
rect 540 637 560 657
rect 580 637 600 657
rect 620 637 640 657
rect 660 637 680 657
rect 700 637 720 657
rect 740 637 760 657
rect 780 637 800 657
rect 820 637 840 657
rect 860 637 880 657
rect 900 637 920 657
rect 940 637 960 657
rect 980 637 1000 657
rect 1020 637 1040 657
rect 1060 637 1080 657
rect 1100 637 1120 657
rect 1140 637 1160 657
rect 1180 637 1200 657
rect 1220 637 1240 657
rect 1260 637 1280 657
rect 1300 637 1320 657
rect 1340 637 1360 657
rect 1380 637 1400 657
rect 1420 637 1440 657
rect 1460 637 1480 657
rect 1500 637 1520 657
rect 1540 637 1560 657
rect 1580 637 1600 657
rect 1620 637 1640 657
rect 1660 637 1680 657
rect 1700 637 1720 657
rect 1740 637 1760 657
rect 1780 637 1800 657
rect 1820 637 1840 657
rect 1860 637 1880 657
rect 1900 637 1920 657
rect 1940 637 1960 657
rect 1980 637 2000 657
rect 2020 637 2040 657
rect 2060 637 2080 657
rect 2100 637 2120 657
rect 2140 637 2160 657
rect 2180 637 2200 657
rect 2220 637 2240 657
rect 2260 637 2280 657
rect 2300 637 2320 657
rect 2340 637 2360 657
rect 2380 637 2400 657
rect 2420 637 2440 657
rect 2460 637 2480 657
rect 2500 637 2520 657
rect 2540 637 2560 657
rect 2580 637 2600 657
rect 2620 637 2640 657
rect 2660 637 2675 657
rect 175 627 2675 637
rect 0 615 155 625
rect 0 595 10 615
rect 30 595 50 615
rect 70 595 90 615
rect 110 595 130 615
rect 0 585 155 595
rect 175 575 2675 585
rect 175 555 200 575
rect 220 555 240 575
rect 260 555 280 575
rect 300 555 320 575
rect 340 555 360 575
rect 380 555 400 575
rect 420 555 440 575
rect 460 555 480 575
rect 500 555 520 575
rect 540 555 560 575
rect 580 555 600 575
rect 620 555 640 575
rect 660 555 680 575
rect 700 555 720 575
rect 740 555 760 575
rect 780 555 800 575
rect 820 555 840 575
rect 860 555 880 575
rect 900 555 920 575
rect 940 555 960 575
rect 980 555 1000 575
rect 1020 555 1040 575
rect 1060 555 1080 575
rect 1100 555 1120 575
rect 1140 555 1160 575
rect 1180 555 1200 575
rect 1220 555 1240 575
rect 1260 555 1280 575
rect 1300 555 1320 575
rect 1340 555 1360 575
rect 1380 555 1400 575
rect 1420 555 1440 575
rect 1460 555 1480 575
rect 1500 555 1520 575
rect 1540 555 1560 575
rect 1580 555 1600 575
rect 1620 555 1640 575
rect 1660 555 1680 575
rect 1700 555 1720 575
rect 1740 555 1760 575
rect 1780 555 1800 575
rect 1820 555 1840 575
rect 1860 555 1880 575
rect 1900 555 1920 575
rect 1940 555 1960 575
rect 1980 555 2000 575
rect 2020 555 2040 575
rect 2060 555 2080 575
rect 2100 555 2120 575
rect 2140 555 2160 575
rect 2180 555 2200 575
rect 2220 555 2240 575
rect 2260 555 2280 575
rect 2300 555 2320 575
rect 2340 555 2360 575
rect 2380 555 2400 575
rect 2420 555 2440 575
rect 2460 555 2480 575
rect 2500 555 2520 575
rect 2540 555 2560 575
rect 2580 555 2600 575
rect 2620 555 2640 575
rect 2660 555 2675 575
rect 175 545 2675 555
rect 0 535 155 545
rect 0 515 10 535
rect 30 515 50 535
rect 70 515 90 535
rect 110 515 130 535
rect 0 505 155 515
rect 175 493 2675 503
rect 175 473 200 493
rect 220 473 240 493
rect 260 473 280 493
rect 300 473 320 493
rect 340 473 360 493
rect 380 473 400 493
rect 420 473 440 493
rect 460 473 480 493
rect 500 473 520 493
rect 540 473 560 493
rect 580 473 600 493
rect 620 473 640 493
rect 660 473 680 493
rect 700 473 720 493
rect 740 473 760 493
rect 780 473 800 493
rect 820 473 840 493
rect 860 473 880 493
rect 900 473 920 493
rect 940 473 960 493
rect 980 473 1000 493
rect 1020 473 1040 493
rect 1060 473 1080 493
rect 1100 473 1120 493
rect 1140 473 1160 493
rect 1180 473 1200 493
rect 1220 473 1240 493
rect 1260 473 1280 493
rect 1300 473 1320 493
rect 1340 473 1360 493
rect 1380 473 1400 493
rect 1420 473 1440 493
rect 1460 473 1480 493
rect 1500 473 1520 493
rect 1540 473 1560 493
rect 1580 473 1600 493
rect 1620 473 1640 493
rect 1660 473 1680 493
rect 1700 473 1720 493
rect 1740 473 1760 493
rect 1780 473 1800 493
rect 1820 473 1840 493
rect 1860 473 1880 493
rect 1900 473 1920 493
rect 1940 473 1960 493
rect 1980 473 2000 493
rect 2020 473 2040 493
rect 2060 473 2080 493
rect 2100 473 2120 493
rect 2140 473 2160 493
rect 2180 473 2200 493
rect 2220 473 2240 493
rect 2260 473 2280 493
rect 2300 473 2320 493
rect 2340 473 2360 493
rect 2380 473 2400 493
rect 2420 473 2440 493
rect 2460 473 2480 493
rect 2500 473 2520 493
rect 2540 473 2560 493
rect 2580 473 2600 493
rect 2620 473 2640 493
rect 2660 473 2675 493
rect 0 455 155 465
rect 175 463 2675 473
rect 0 435 10 455
rect 30 435 50 455
rect 70 435 90 455
rect 110 435 130 455
rect 0 425 155 435
rect 175 411 2675 421
rect 175 391 200 411
rect 220 391 240 411
rect 260 391 280 411
rect 300 391 320 411
rect 340 391 360 411
rect 380 391 400 411
rect 420 391 440 411
rect 460 391 480 411
rect 500 391 520 411
rect 540 391 560 411
rect 580 391 600 411
rect 620 391 640 411
rect 660 391 680 411
rect 700 391 720 411
rect 740 391 760 411
rect 780 391 800 411
rect 820 391 840 411
rect 860 391 880 411
rect 900 391 920 411
rect 940 391 960 411
rect 980 391 1000 411
rect 1020 391 1040 411
rect 1060 391 1080 411
rect 1100 391 1120 411
rect 1140 391 1160 411
rect 1180 391 1200 411
rect 1220 391 1240 411
rect 1260 391 1280 411
rect 1300 391 1320 411
rect 1340 391 1360 411
rect 1380 391 1400 411
rect 1420 391 1440 411
rect 1460 391 1480 411
rect 1500 391 1520 411
rect 1540 391 1560 411
rect 1580 391 1600 411
rect 1620 391 1640 411
rect 1660 391 1680 411
rect 1700 391 1720 411
rect 1740 391 1760 411
rect 1780 391 1800 411
rect 1820 391 1840 411
rect 1860 391 1880 411
rect 1900 391 1920 411
rect 1940 391 1960 411
rect 1980 391 2000 411
rect 2020 391 2040 411
rect 2060 391 2080 411
rect 2100 391 2120 411
rect 2140 391 2160 411
rect 2180 391 2200 411
rect 2220 391 2240 411
rect 2260 391 2280 411
rect 2300 391 2320 411
rect 2340 391 2360 411
rect 2380 391 2400 411
rect 2420 391 2440 411
rect 2460 391 2480 411
rect 2500 391 2520 411
rect 2540 391 2560 411
rect 2580 391 2600 411
rect 2620 391 2640 411
rect 2660 391 2675 411
rect 175 381 2675 391
rect 0 370 155 380
rect 0 350 10 370
rect 30 350 50 370
rect 70 350 90 370
rect 110 350 130 370
rect 0 340 155 350
rect 175 329 2675 339
rect 175 309 200 329
rect 220 309 240 329
rect 260 309 280 329
rect 300 309 320 329
rect 340 309 360 329
rect 380 309 400 329
rect 420 309 440 329
rect 460 309 480 329
rect 500 309 520 329
rect 540 309 560 329
rect 580 309 600 329
rect 620 309 640 329
rect 660 309 680 329
rect 700 309 720 329
rect 740 309 760 329
rect 780 309 800 329
rect 820 309 840 329
rect 860 309 880 329
rect 900 309 920 329
rect 940 309 960 329
rect 980 309 1000 329
rect 1020 309 1040 329
rect 1060 309 1080 329
rect 1100 309 1120 329
rect 1140 309 1160 329
rect 1180 309 1200 329
rect 1220 309 1240 329
rect 1260 309 1280 329
rect 1300 309 1320 329
rect 1340 309 1360 329
rect 1380 309 1400 329
rect 1420 309 1440 329
rect 1460 309 1480 329
rect 1500 309 1520 329
rect 1540 309 1560 329
rect 1580 309 1600 329
rect 1620 309 1640 329
rect 1660 309 1680 329
rect 1700 309 1720 329
rect 1740 309 1760 329
rect 1780 309 1800 329
rect 1820 309 1840 329
rect 1860 309 1880 329
rect 1900 309 1920 329
rect 1940 309 1960 329
rect 1980 309 2000 329
rect 2020 309 2040 329
rect 2060 309 2080 329
rect 2100 309 2120 329
rect 2140 309 2160 329
rect 2180 309 2200 329
rect 2220 309 2240 329
rect 2260 309 2280 329
rect 2300 309 2320 329
rect 2340 309 2360 329
rect 2380 309 2400 329
rect 2420 309 2440 329
rect 2460 309 2480 329
rect 2500 309 2520 329
rect 2540 309 2560 329
rect 2580 309 2600 329
rect 2620 309 2640 329
rect 2660 309 2675 329
rect 0 290 155 300
rect 175 299 2675 309
rect 0 270 10 290
rect 30 270 50 290
rect 70 270 90 290
rect 110 270 130 290
rect 0 260 155 270
rect 175 247 2675 257
rect 175 227 200 247
rect 220 227 240 247
rect 260 227 280 247
rect 300 227 320 247
rect 340 227 360 247
rect 380 227 400 247
rect 420 227 440 247
rect 460 227 480 247
rect 500 227 520 247
rect 540 227 560 247
rect 580 227 600 247
rect 620 227 640 247
rect 660 227 680 247
rect 700 227 720 247
rect 740 227 760 247
rect 780 227 800 247
rect 820 227 840 247
rect 860 227 880 247
rect 900 227 920 247
rect 940 227 960 247
rect 980 227 1000 247
rect 1020 227 1040 247
rect 1060 227 1080 247
rect 1100 227 1120 247
rect 1140 227 1160 247
rect 1180 227 1200 247
rect 1220 227 1240 247
rect 1260 227 1280 247
rect 1300 227 1320 247
rect 1340 227 1360 247
rect 1380 227 1400 247
rect 1420 227 1440 247
rect 1460 227 1480 247
rect 1500 227 1520 247
rect 1540 227 1560 247
rect 1580 227 1600 247
rect 1620 227 1640 247
rect 1660 227 1680 247
rect 1700 227 1720 247
rect 1740 227 1760 247
rect 1780 227 1800 247
rect 1820 227 1840 247
rect 1860 227 1880 247
rect 1900 227 1920 247
rect 1940 227 1960 247
rect 1980 227 2000 247
rect 2020 227 2040 247
rect 2060 227 2080 247
rect 2100 227 2120 247
rect 2140 227 2160 247
rect 2180 227 2200 247
rect 2220 227 2240 247
rect 2260 227 2280 247
rect 2300 227 2320 247
rect 2340 227 2360 247
rect 2380 227 2400 247
rect 2420 227 2440 247
rect 2460 227 2480 247
rect 2500 227 2520 247
rect 2540 227 2560 247
rect 2580 227 2600 247
rect 2620 227 2640 247
rect 2660 227 2675 247
rect 0 210 155 220
rect 175 217 2675 227
rect 0 190 10 210
rect 30 190 50 210
rect 70 190 90 210
rect 110 190 130 210
rect 0 180 155 190
rect 175 165 2675 175
rect 175 145 200 165
rect 220 145 240 165
rect 260 145 280 165
rect 300 145 320 165
rect 340 145 360 165
rect 380 145 400 165
rect 420 145 440 165
rect 460 145 480 165
rect 500 145 520 165
rect 540 145 560 165
rect 580 145 600 165
rect 620 145 640 165
rect 660 145 680 165
rect 700 145 720 165
rect 740 145 760 165
rect 780 145 800 165
rect 820 145 840 165
rect 860 145 880 165
rect 900 145 920 165
rect 940 145 960 165
rect 980 145 1000 165
rect 1020 145 1040 165
rect 1060 145 1080 165
rect 1100 145 1120 165
rect 1140 145 1160 165
rect 1180 145 1200 165
rect 1220 145 1240 165
rect 1260 145 1280 165
rect 1300 145 1320 165
rect 1340 145 1360 165
rect 1380 145 1400 165
rect 1420 145 1440 165
rect 1460 145 1480 165
rect 1500 145 1520 165
rect 1540 145 1560 165
rect 1580 145 1600 165
rect 1620 145 1640 165
rect 1660 145 1680 165
rect 1700 145 1720 165
rect 1740 145 1760 165
rect 1780 145 1800 165
rect 1820 145 1840 165
rect 1860 145 1880 165
rect 1900 145 1920 165
rect 1940 145 1960 165
rect 1980 145 2000 165
rect 2020 145 2040 165
rect 2060 145 2080 165
rect 2100 145 2120 165
rect 2140 145 2160 165
rect 2180 145 2200 165
rect 2220 145 2240 165
rect 2260 145 2280 165
rect 2300 145 2320 165
rect 2340 145 2360 165
rect 2380 145 2400 165
rect 2420 145 2440 165
rect 2460 145 2480 165
rect 2500 145 2520 165
rect 2540 145 2560 165
rect 2580 145 2600 165
rect 2620 145 2640 165
rect 2660 145 2675 165
rect 175 135 2675 145
rect 175 95 2675 105
rect 175 75 200 95
rect 220 75 240 95
rect 260 75 280 95
rect 300 75 320 95
rect 340 75 360 95
rect 380 75 400 95
rect 420 75 440 95
rect 460 75 480 95
rect 500 75 520 95
rect 540 75 560 95
rect 580 75 600 95
rect 620 75 640 95
rect 660 75 680 95
rect 700 75 720 95
rect 740 75 760 95
rect 780 75 800 95
rect 820 75 840 95
rect 860 75 880 95
rect 900 75 920 95
rect 940 75 960 95
rect 980 75 1000 95
rect 1020 75 1040 95
rect 1060 75 1080 95
rect 1100 75 1120 95
rect 1140 75 1160 95
rect 1180 75 1200 95
rect 1220 75 1240 95
rect 1260 75 1280 95
rect 1300 75 1320 95
rect 1340 75 1360 95
rect 1380 75 1400 95
rect 1420 75 1440 95
rect 1460 75 1480 95
rect 1500 75 1520 95
rect 1540 75 1560 95
rect 1580 75 1600 95
rect 1620 75 1640 95
rect 1660 75 1680 95
rect 1700 75 1720 95
rect 1740 75 1760 95
rect 1780 75 1800 95
rect 1820 75 1840 95
rect 1860 75 1880 95
rect 1900 75 1920 95
rect 1940 75 1960 95
rect 1980 75 2000 95
rect 2020 75 2040 95
rect 2060 75 2080 95
rect 2100 75 2120 95
rect 2140 75 2160 95
rect 2180 75 2200 95
rect 2220 75 2240 95
rect 2260 75 2280 95
rect 2300 75 2320 95
rect 2340 75 2360 95
rect 2380 75 2400 95
rect 2420 75 2440 95
rect 2460 75 2480 95
rect 2500 75 2520 95
rect 2540 75 2560 95
rect 2580 75 2600 95
rect 2620 75 2640 95
rect 2660 75 2675 95
rect 175 65 2675 75
rect 105 -10 2605 0
rect 105 -30 120 -10
rect 140 -30 160 -10
rect 180 -30 200 -10
rect 220 -30 240 -10
rect 260 -30 280 -10
rect 300 -30 320 -10
rect 340 -30 360 -10
rect 380 -30 400 -10
rect 420 -30 440 -10
rect 460 -30 480 -10
rect 500 -30 520 -10
rect 540 -30 560 -10
rect 580 -30 600 -10
rect 620 -30 640 -10
rect 660 -30 680 -10
rect 700 -30 720 -10
rect 740 -30 760 -10
rect 780 -30 800 -10
rect 820 -30 840 -10
rect 860 -30 880 -10
rect 900 -30 920 -10
rect 940 -30 960 -10
rect 980 -30 1000 -10
rect 1020 -30 1040 -10
rect 1060 -30 1080 -10
rect 1100 -30 1120 -10
rect 1140 -30 1160 -10
rect 1180 -30 1200 -10
rect 1220 -30 1240 -10
rect 1260 -30 1280 -10
rect 1300 -30 1320 -10
rect 1340 -30 1360 -10
rect 1380 -30 1400 -10
rect 1420 -30 1440 -10
rect 1460 -30 1480 -10
rect 1500 -30 1520 -10
rect 1540 -30 1560 -10
rect 1580 -30 1600 -10
rect 1620 -30 1640 -10
rect 1660 -30 1680 -10
rect 1700 -30 1720 -10
rect 1740 -30 1760 -10
rect 1780 -30 1800 -10
rect 1820 -30 1840 -10
rect 1860 -30 1880 -10
rect 1900 -30 1920 -10
rect 1940 -30 1960 -10
rect 1980 -30 2000 -10
rect 2020 -30 2040 -10
rect 2060 -30 2080 -10
rect 2100 -30 2120 -10
rect 2140 -30 2160 -10
rect 2180 -30 2200 -10
rect 2220 -30 2240 -10
rect 2260 -30 2280 -10
rect 2300 -30 2320 -10
rect 2340 -30 2360 -10
rect 2380 -30 2400 -10
rect 2420 -30 2440 -10
rect 2460 -30 2480 -10
rect 2500 -30 2520 -10
rect 2540 -30 2560 -10
rect 2590 -30 2605 -10
rect 105 -50 2605 -30
rect 105 -70 120 -50
rect 140 -70 160 -50
rect 180 -70 200 -50
rect 220 -70 240 -50
rect 260 -70 280 -50
rect 300 -70 320 -50
rect 340 -70 360 -50
rect 380 -70 400 -50
rect 420 -70 440 -50
rect 460 -70 480 -50
rect 500 -70 520 -50
rect 540 -70 560 -50
rect 580 -70 600 -50
rect 620 -70 640 -50
rect 660 -70 680 -50
rect 700 -70 720 -50
rect 740 -70 760 -50
rect 780 -70 800 -50
rect 820 -70 840 -50
rect 860 -70 880 -50
rect 900 -70 920 -50
rect 940 -70 960 -50
rect 980 -70 1000 -50
rect 1020 -70 1040 -50
rect 1060 -70 1080 -50
rect 1100 -70 1120 -50
rect 1140 -70 1160 -50
rect 1180 -70 1200 -50
rect 1220 -70 1240 -50
rect 1260 -70 1280 -50
rect 1300 -70 1320 -50
rect 1340 -70 1360 -50
rect 1380 -70 1400 -50
rect 1420 -70 1440 -50
rect 1460 -70 1480 -50
rect 1500 -70 1520 -50
rect 1540 -70 1560 -50
rect 1580 -70 1600 -50
rect 1620 -70 1640 -50
rect 1660 -70 1680 -50
rect 1700 -70 1720 -50
rect 1740 -70 1760 -50
rect 1780 -70 1800 -50
rect 1820 -70 1840 -50
rect 1860 -70 1880 -50
rect 1900 -70 1920 -50
rect 1940 -70 1960 -50
rect 1980 -70 2000 -50
rect 2020 -70 2040 -50
rect 2060 -70 2080 -50
rect 2100 -70 2120 -50
rect 2140 -70 2160 -50
rect 2180 -70 2200 -50
rect 2220 -70 2240 -50
rect 2260 -70 2280 -50
rect 2300 -70 2320 -50
rect 2340 -70 2360 -50
rect 2380 -70 2400 -50
rect 2420 -70 2440 -50
rect 2460 -70 2480 -50
rect 2500 -70 2520 -50
rect 2540 -70 2560 -50
rect 2590 -70 2605 -50
rect 105 -80 2605 -70
rect -70 -95 85 -85
rect -70 -120 -60 -95
rect -40 -120 -20 -95
rect 0 -120 20 -95
rect 40 -120 60 -95
rect -70 -130 85 -120
rect 105 -145 2605 -135
rect 105 -165 120 -145
rect 140 -165 160 -145
rect 180 -165 200 -145
rect 220 -165 240 -145
rect 260 -165 280 -145
rect 300 -165 320 -145
rect 340 -165 360 -145
rect 380 -165 400 -145
rect 420 -165 440 -145
rect 460 -165 480 -145
rect 500 -165 520 -145
rect 540 -165 560 -145
rect 580 -165 600 -145
rect 620 -165 640 -145
rect 660 -165 680 -145
rect 700 -165 720 -145
rect 740 -165 760 -145
rect 780 -165 800 -145
rect 820 -165 840 -145
rect 860 -165 880 -145
rect 900 -165 920 -145
rect 940 -165 960 -145
rect 980 -165 1000 -145
rect 1020 -165 1040 -145
rect 1060 -165 1080 -145
rect 1100 -165 1120 -145
rect 1140 -165 1160 -145
rect 1180 -165 1200 -145
rect 1220 -165 1240 -145
rect 1260 -165 1280 -145
rect 1300 -165 1320 -145
rect 1340 -165 1360 -145
rect 1380 -165 1400 -145
rect 1420 -165 1440 -145
rect 1460 -165 1480 -145
rect 1500 -165 1520 -145
rect 1540 -165 1560 -145
rect 1580 -165 1600 -145
rect 1620 -165 1640 -145
rect 1660 -165 1680 -145
rect 1700 -165 1720 -145
rect 1740 -165 1760 -145
rect 1780 -165 1800 -145
rect 1820 -165 1840 -145
rect 1860 -165 1880 -145
rect 1900 -165 1920 -145
rect 1940 -165 1960 -145
rect 1980 -165 2000 -145
rect 2020 -165 2040 -145
rect 2060 -165 2080 -145
rect 2100 -165 2120 -145
rect 2140 -165 2160 -145
rect 2180 -165 2200 -145
rect 2220 -165 2240 -145
rect 2260 -165 2280 -145
rect 2300 -165 2320 -145
rect 2340 -165 2360 -145
rect 2380 -165 2400 -145
rect 2420 -165 2440 -145
rect 2460 -165 2480 -145
rect 2500 -165 2520 -145
rect 2540 -165 2560 -145
rect 2590 -165 2605 -145
rect 105 -175 2605 -165
rect -70 -190 85 -180
rect -70 -215 -60 -190
rect -40 -215 -20 -190
rect 0 -215 20 -190
rect 40 -215 60 -190
rect -70 -225 85 -215
rect 105 -240 2605 -230
rect 105 -260 120 -240
rect 140 -260 160 -240
rect 180 -260 200 -240
rect 220 -260 240 -240
rect 260 -260 280 -240
rect 300 -260 320 -240
rect 340 -260 360 -240
rect 380 -260 400 -240
rect 420 -260 440 -240
rect 460 -260 480 -240
rect 500 -260 520 -240
rect 540 -260 560 -240
rect 580 -260 600 -240
rect 620 -260 640 -240
rect 660 -260 680 -240
rect 700 -260 720 -240
rect 740 -260 760 -240
rect 780 -260 800 -240
rect 820 -260 840 -240
rect 860 -260 880 -240
rect 900 -260 920 -240
rect 940 -260 960 -240
rect 980 -260 1000 -240
rect 1020 -260 1040 -240
rect 1060 -260 1080 -240
rect 1100 -260 1120 -240
rect 1140 -260 1160 -240
rect 1180 -260 1200 -240
rect 1220 -260 1240 -240
rect 1260 -260 1280 -240
rect 1300 -260 1320 -240
rect 1340 -260 1360 -240
rect 1380 -260 1400 -240
rect 1420 -260 1440 -240
rect 1460 -260 1480 -240
rect 1500 -260 1520 -240
rect 1540 -260 1560 -240
rect 1580 -260 1600 -240
rect 1620 -260 1640 -240
rect 1660 -260 1680 -240
rect 1700 -260 1720 -240
rect 1740 -260 1760 -240
rect 1780 -260 1800 -240
rect 1820 -260 1840 -240
rect 1860 -260 1880 -240
rect 1900 -260 1920 -240
rect 1940 -260 1960 -240
rect 1980 -260 2000 -240
rect 2020 -260 2040 -240
rect 2060 -260 2080 -240
rect 2100 -260 2120 -240
rect 2140 -260 2160 -240
rect 2180 -260 2200 -240
rect 2220 -260 2240 -240
rect 2260 -260 2280 -240
rect 2300 -260 2320 -240
rect 2340 -260 2360 -240
rect 2380 -260 2400 -240
rect 2420 -260 2440 -240
rect 2460 -260 2480 -240
rect 2500 -260 2520 -240
rect 2540 -260 2560 -240
rect 2590 -260 2605 -240
rect 105 -270 2605 -260
rect -70 -285 85 -275
rect -70 -310 -60 -285
rect -40 -310 -20 -285
rect 0 -310 20 -285
rect 40 -310 60 -285
rect -70 -320 85 -310
rect 105 -335 2605 -325
rect 105 -355 120 -335
rect 140 -355 160 -335
rect 180 -355 200 -335
rect 220 -355 240 -335
rect 260 -355 280 -335
rect 300 -355 320 -335
rect 340 -355 360 -335
rect 380 -355 400 -335
rect 420 -355 440 -335
rect 460 -355 480 -335
rect 500 -355 520 -335
rect 540 -355 560 -335
rect 580 -355 600 -335
rect 620 -355 640 -335
rect 660 -355 680 -335
rect 700 -355 720 -335
rect 740 -355 760 -335
rect 780 -355 800 -335
rect 820 -355 840 -335
rect 860 -355 880 -335
rect 900 -355 920 -335
rect 940 -355 960 -335
rect 980 -355 1000 -335
rect 1020 -355 1040 -335
rect 1060 -355 1080 -335
rect 1100 -355 1120 -335
rect 1140 -355 1160 -335
rect 1180 -355 1200 -335
rect 1220 -355 1240 -335
rect 1260 -355 1280 -335
rect 1300 -355 1320 -335
rect 1340 -355 1360 -335
rect 1380 -355 1400 -335
rect 1420 -355 1440 -335
rect 1460 -355 1480 -335
rect 1500 -355 1520 -335
rect 1540 -355 1560 -335
rect 1580 -355 1600 -335
rect 1620 -355 1640 -335
rect 1660 -355 1680 -335
rect 1700 -355 1720 -335
rect 1740 -355 1760 -335
rect 1780 -355 1800 -335
rect 1820 -355 1840 -335
rect 1860 -355 1880 -335
rect 1900 -355 1920 -335
rect 1940 -355 1960 -335
rect 1980 -355 2000 -335
rect 2020 -355 2040 -335
rect 2060 -355 2080 -335
rect 2100 -355 2120 -335
rect 2140 -355 2160 -335
rect 2180 -355 2200 -335
rect 2220 -355 2240 -335
rect 2260 -355 2280 -335
rect 2300 -355 2320 -335
rect 2340 -355 2360 -335
rect 2380 -355 2400 -335
rect 2420 -355 2440 -335
rect 2460 -355 2480 -335
rect 2500 -355 2520 -335
rect 2540 -355 2560 -335
rect 2590 -355 2605 -335
rect 105 -365 2605 -355
rect -70 -380 85 -370
rect -70 -405 -60 -380
rect -40 -405 -20 -380
rect 0 -405 20 -380
rect 40 -405 60 -380
rect -70 -415 85 -405
rect 105 -430 2605 -420
rect 105 -450 120 -430
rect 140 -450 160 -430
rect 180 -450 200 -430
rect 220 -450 240 -430
rect 260 -450 280 -430
rect 300 -450 320 -430
rect 340 -450 360 -430
rect 380 -450 400 -430
rect 420 -450 440 -430
rect 460 -450 480 -430
rect 500 -450 520 -430
rect 540 -450 560 -430
rect 580 -450 600 -430
rect 620 -450 640 -430
rect 660 -450 680 -430
rect 700 -450 720 -430
rect 740 -450 760 -430
rect 780 -450 800 -430
rect 820 -450 840 -430
rect 860 -450 880 -430
rect 900 -450 920 -430
rect 940 -450 960 -430
rect 980 -450 1000 -430
rect 1020 -450 1040 -430
rect 1060 -450 1080 -430
rect 1100 -450 1120 -430
rect 1140 -450 1160 -430
rect 1180 -450 1200 -430
rect 1220 -450 1240 -430
rect 1260 -450 1280 -430
rect 1300 -450 1320 -430
rect 1340 -450 1360 -430
rect 1380 -450 1400 -430
rect 1420 -450 1440 -430
rect 1460 -450 1480 -430
rect 1500 -450 1520 -430
rect 1540 -450 1560 -430
rect 1580 -450 1600 -430
rect 1620 -450 1640 -430
rect 1660 -450 1680 -430
rect 1700 -450 1720 -430
rect 1740 -450 1760 -430
rect 1780 -450 1800 -430
rect 1820 -450 1840 -430
rect 1860 -450 1880 -430
rect 1900 -450 1920 -430
rect 1940 -450 1960 -430
rect 1980 -450 2000 -430
rect 2020 -450 2040 -430
rect 2060 -450 2080 -430
rect 2100 -450 2120 -430
rect 2140 -450 2160 -430
rect 2180 -450 2200 -430
rect 2220 -450 2240 -430
rect 2260 -450 2280 -430
rect 2300 -450 2320 -430
rect 2340 -450 2360 -430
rect 2380 -450 2400 -430
rect 2420 -450 2440 -430
rect 2460 -450 2480 -430
rect 2500 -450 2520 -430
rect 2540 -450 2560 -430
rect 2590 -450 2605 -430
rect 105 -460 2605 -450
rect -70 -475 85 -465
rect -70 -500 -60 -475
rect -40 -500 -20 -475
rect 0 -500 20 -475
rect 40 -500 60 -475
rect -70 -510 85 -500
rect 105 -525 2605 -515
rect 105 -545 120 -525
rect 140 -545 160 -525
rect 180 -545 200 -525
rect 220 -545 240 -525
rect 260 -545 280 -525
rect 300 -545 320 -525
rect 340 -545 360 -525
rect 380 -545 400 -525
rect 420 -545 440 -525
rect 460 -545 480 -525
rect 500 -545 520 -525
rect 540 -545 560 -525
rect 580 -545 600 -525
rect 620 -545 640 -525
rect 660 -545 680 -525
rect 700 -545 720 -525
rect 740 -545 760 -525
rect 780 -545 800 -525
rect 820 -545 840 -525
rect 860 -545 880 -525
rect 900 -545 920 -525
rect 940 -545 960 -525
rect 980 -545 1000 -525
rect 1020 -545 1040 -525
rect 1060 -545 1080 -525
rect 1100 -545 1120 -525
rect 1140 -545 1160 -525
rect 1180 -545 1200 -525
rect 1220 -545 1240 -525
rect 1260 -545 1280 -525
rect 1300 -545 1320 -525
rect 1340 -545 1360 -525
rect 1380 -545 1400 -525
rect 1420 -545 1440 -525
rect 1460 -545 1480 -525
rect 1500 -545 1520 -525
rect 1540 -545 1560 -525
rect 1580 -545 1600 -525
rect 1620 -545 1640 -525
rect 1660 -545 1680 -525
rect 1700 -545 1720 -525
rect 1740 -545 1760 -525
rect 1780 -545 1800 -525
rect 1820 -545 1840 -525
rect 1860 -545 1880 -525
rect 1900 -545 1920 -525
rect 1940 -545 1960 -525
rect 1980 -545 2000 -525
rect 2020 -545 2040 -525
rect 2060 -545 2080 -525
rect 2100 -545 2120 -525
rect 2140 -545 2160 -525
rect 2180 -545 2200 -525
rect 2220 -545 2240 -525
rect 2260 -545 2280 -525
rect 2300 -545 2320 -525
rect 2340 -545 2360 -525
rect 2380 -545 2400 -525
rect 2420 -545 2440 -525
rect 2460 -545 2480 -525
rect 2500 -545 2520 -525
rect 2540 -545 2560 -525
rect 2590 -545 2605 -525
rect 105 -555 2605 -545
rect -70 -570 85 -560
rect -70 -595 -60 -570
rect -40 -595 -20 -570
rect 0 -595 20 -570
rect 40 -595 60 -570
rect -70 -605 85 -595
rect 105 -620 2605 -610
rect 105 -640 120 -620
rect 140 -640 160 -620
rect 180 -640 200 -620
rect 220 -640 240 -620
rect 260 -640 280 -620
rect 300 -640 320 -620
rect 340 -640 360 -620
rect 380 -640 400 -620
rect 420 -640 440 -620
rect 460 -640 480 -620
rect 500 -640 520 -620
rect 540 -640 560 -620
rect 580 -640 600 -620
rect 620 -640 640 -620
rect 660 -640 680 -620
rect 700 -640 720 -620
rect 740 -640 760 -620
rect 780 -640 800 -620
rect 820 -640 840 -620
rect 860 -640 880 -620
rect 900 -640 920 -620
rect 940 -640 960 -620
rect 980 -640 1000 -620
rect 1020 -640 1040 -620
rect 1060 -640 1080 -620
rect 1100 -640 1120 -620
rect 1140 -640 1160 -620
rect 1180 -640 1200 -620
rect 1220 -640 1240 -620
rect 1260 -640 1280 -620
rect 1300 -640 1320 -620
rect 1340 -640 1360 -620
rect 1380 -640 1400 -620
rect 1420 -640 1440 -620
rect 1460 -640 1480 -620
rect 1500 -640 1520 -620
rect 1540 -640 1560 -620
rect 1580 -640 1600 -620
rect 1620 -640 1640 -620
rect 1660 -640 1680 -620
rect 1700 -640 1720 -620
rect 1740 -640 1760 -620
rect 1780 -640 1800 -620
rect 1820 -640 1840 -620
rect 1860 -640 1880 -620
rect 1900 -640 1920 -620
rect 1940 -640 1960 -620
rect 1980 -640 2000 -620
rect 2020 -640 2040 -620
rect 2060 -640 2080 -620
rect 2100 -640 2120 -620
rect 2140 -640 2160 -620
rect 2180 -640 2200 -620
rect 2220 -640 2240 -620
rect 2260 -640 2280 -620
rect 2300 -640 2320 -620
rect 2340 -640 2360 -620
rect 2380 -640 2400 -620
rect 2420 -640 2440 -620
rect 2460 -640 2480 -620
rect 2500 -640 2520 -620
rect 2540 -640 2560 -620
rect 2590 -640 2605 -620
rect 105 -650 2605 -640
rect -70 -665 85 -655
rect -70 -690 -60 -665
rect -40 -690 -20 -665
rect 0 -690 20 -665
rect 40 -690 60 -665
rect -70 -700 85 -690
rect 105 -715 2605 -705
rect 105 -735 120 -715
rect 140 -735 160 -715
rect 180 -735 200 -715
rect 220 -735 240 -715
rect 260 -735 280 -715
rect 300 -735 320 -715
rect 340 -735 360 -715
rect 380 -735 400 -715
rect 420 -735 440 -715
rect 460 -735 480 -715
rect 500 -735 520 -715
rect 540 -735 560 -715
rect 580 -735 600 -715
rect 620 -735 640 -715
rect 660 -735 680 -715
rect 700 -735 720 -715
rect 740 -735 760 -715
rect 780 -735 800 -715
rect 820 -735 840 -715
rect 860 -735 880 -715
rect 900 -735 920 -715
rect 940 -735 960 -715
rect 980 -735 1000 -715
rect 1020 -735 1040 -715
rect 1060 -735 1080 -715
rect 1100 -735 1120 -715
rect 1140 -735 1160 -715
rect 1180 -735 1200 -715
rect 1220 -735 1240 -715
rect 1260 -735 1280 -715
rect 1300 -735 1320 -715
rect 1340 -735 1360 -715
rect 1380 -735 1400 -715
rect 1420 -735 1440 -715
rect 1460 -735 1480 -715
rect 1500 -735 1520 -715
rect 1540 -735 1560 -715
rect 1580 -735 1600 -715
rect 1620 -735 1640 -715
rect 1660 -735 1680 -715
rect 1700 -735 1720 -715
rect 1740 -735 1760 -715
rect 1780 -735 1800 -715
rect 1820 -735 1840 -715
rect 1860 -735 1880 -715
rect 1900 -735 1920 -715
rect 1940 -735 1960 -715
rect 1980 -735 2000 -715
rect 2020 -735 2040 -715
rect 2060 -735 2080 -715
rect 2100 -735 2120 -715
rect 2140 -735 2160 -715
rect 2180 -735 2200 -715
rect 2220 -735 2240 -715
rect 2260 -735 2280 -715
rect 2300 -735 2320 -715
rect 2340 -735 2360 -715
rect 2380 -735 2400 -715
rect 2420 -735 2440 -715
rect 2460 -735 2480 -715
rect 2500 -735 2520 -715
rect 2540 -735 2560 -715
rect 2590 -735 2605 -715
rect 105 -745 2605 -735
rect -70 -760 85 -750
rect -70 -785 -60 -760
rect -40 -785 -20 -760
rect 0 -785 20 -760
rect 40 -785 60 -760
rect -70 -795 85 -785
rect 105 -810 2605 -800
rect 105 -830 120 -810
rect 140 -830 160 -810
rect 180 -830 200 -810
rect 220 -830 240 -810
rect 260 -830 280 -810
rect 300 -830 320 -810
rect 340 -830 360 -810
rect 380 -830 400 -810
rect 420 -830 440 -810
rect 460 -830 480 -810
rect 500 -830 520 -810
rect 540 -830 560 -810
rect 580 -830 600 -810
rect 620 -830 640 -810
rect 660 -830 680 -810
rect 700 -830 720 -810
rect 740 -830 760 -810
rect 780 -830 800 -810
rect 820 -830 840 -810
rect 860 -830 880 -810
rect 900 -830 920 -810
rect 940 -830 960 -810
rect 980 -830 1000 -810
rect 1020 -830 1040 -810
rect 1060 -830 1080 -810
rect 1100 -830 1120 -810
rect 1140 -830 1160 -810
rect 1180 -830 1200 -810
rect 1220 -830 1240 -810
rect 1260 -830 1280 -810
rect 1300 -830 1320 -810
rect 1340 -830 1360 -810
rect 1380 -830 1400 -810
rect 1420 -830 1440 -810
rect 1460 -830 1480 -810
rect 1500 -830 1520 -810
rect 1540 -830 1560 -810
rect 1580 -830 1600 -810
rect 1620 -830 1640 -810
rect 1660 -830 1680 -810
rect 1700 -830 1720 -810
rect 1740 -830 1760 -810
rect 1780 -830 1800 -810
rect 1820 -830 1840 -810
rect 1860 -830 1880 -810
rect 1900 -830 1920 -810
rect 1940 -830 1960 -810
rect 1980 -830 2000 -810
rect 2020 -830 2040 -810
rect 2060 -830 2080 -810
rect 2100 -830 2120 -810
rect 2140 -830 2160 -810
rect 2180 -830 2200 -810
rect 2220 -830 2240 -810
rect 2260 -830 2280 -810
rect 2300 -830 2320 -810
rect 2340 -830 2360 -810
rect 2380 -830 2400 -810
rect 2420 -830 2440 -810
rect 2460 -830 2480 -810
rect 2500 -830 2520 -810
rect 2540 -830 2560 -810
rect 2590 -830 2605 -810
rect 105 -840 2605 -830
rect -70 -855 85 -845
rect -70 -880 -60 -855
rect -40 -880 -20 -855
rect 0 -880 20 -855
rect 40 -880 60 -855
rect -70 -890 85 -880
rect 105 -905 2605 -895
rect 105 -925 120 -905
rect 140 -925 160 -905
rect 180 -925 200 -905
rect 220 -925 240 -905
rect 260 -925 280 -905
rect 300 -925 320 -905
rect 340 -925 360 -905
rect 380 -925 400 -905
rect 420 -925 440 -905
rect 460 -925 480 -905
rect 500 -925 520 -905
rect 540 -925 560 -905
rect 580 -925 600 -905
rect 620 -925 640 -905
rect 660 -925 680 -905
rect 700 -925 720 -905
rect 740 -925 760 -905
rect 780 -925 800 -905
rect 820 -925 840 -905
rect 860 -925 880 -905
rect 900 -925 920 -905
rect 940 -925 960 -905
rect 980 -925 1000 -905
rect 1020 -925 1040 -905
rect 1060 -925 1080 -905
rect 1100 -925 1120 -905
rect 1140 -925 1160 -905
rect 1180 -925 1200 -905
rect 1220 -925 1240 -905
rect 1260 -925 1280 -905
rect 1300 -925 1320 -905
rect 1340 -925 1360 -905
rect 1380 -925 1400 -905
rect 1420 -925 1440 -905
rect 1460 -925 1480 -905
rect 1500 -925 1520 -905
rect 1540 -925 1560 -905
rect 1580 -925 1600 -905
rect 1620 -925 1640 -905
rect 1660 -925 1680 -905
rect 1700 -925 1720 -905
rect 1740 -925 1760 -905
rect 1780 -925 1800 -905
rect 1820 -925 1840 -905
rect 1860 -925 1880 -905
rect 1900 -925 1920 -905
rect 1940 -925 1960 -905
rect 1980 -925 2000 -905
rect 2020 -925 2040 -905
rect 2060 -925 2080 -905
rect 2100 -925 2120 -905
rect 2140 -925 2160 -905
rect 2180 -925 2200 -905
rect 2220 -925 2240 -905
rect 2260 -925 2280 -905
rect 2300 -925 2320 -905
rect 2340 -925 2360 -905
rect 2380 -925 2400 -905
rect 2420 -925 2440 -905
rect 2460 -925 2480 -905
rect 2500 -925 2520 -905
rect 2540 -925 2560 -905
rect 2590 -925 2605 -905
rect 105 -935 2605 -925
rect -70 -950 85 -940
rect -70 -975 -60 -950
rect -40 -975 -20 -950
rect 0 -975 20 -950
rect 40 -975 60 -950
rect -70 -985 85 -975
rect 105 -1000 2605 -990
rect 105 -1020 120 -1000
rect 140 -1020 160 -1000
rect 180 -1020 200 -1000
rect 220 -1020 240 -1000
rect 260 -1020 280 -1000
rect 300 -1020 320 -1000
rect 340 -1020 360 -1000
rect 380 -1020 400 -1000
rect 420 -1020 440 -1000
rect 460 -1020 480 -1000
rect 500 -1020 520 -1000
rect 540 -1020 560 -1000
rect 580 -1020 600 -1000
rect 620 -1020 640 -1000
rect 660 -1020 680 -1000
rect 700 -1020 720 -1000
rect 740 -1020 760 -1000
rect 780 -1020 800 -1000
rect 820 -1020 840 -1000
rect 860 -1020 880 -1000
rect 900 -1020 920 -1000
rect 940 -1020 960 -1000
rect 980 -1020 1000 -1000
rect 1020 -1020 1040 -1000
rect 1060 -1020 1080 -1000
rect 1100 -1020 1120 -1000
rect 1140 -1020 1160 -1000
rect 1180 -1020 1200 -1000
rect 1220 -1020 1240 -1000
rect 1260 -1020 1280 -1000
rect 1300 -1020 1320 -1000
rect 1340 -1020 1360 -1000
rect 1380 -1020 1400 -1000
rect 1420 -1020 1440 -1000
rect 1460 -1020 1480 -1000
rect 1500 -1020 1520 -1000
rect 1540 -1020 1560 -1000
rect 1580 -1020 1600 -1000
rect 1620 -1020 1640 -1000
rect 1660 -1020 1680 -1000
rect 1700 -1020 1720 -1000
rect 1740 -1020 1760 -1000
rect 1780 -1020 1800 -1000
rect 1820 -1020 1840 -1000
rect 1860 -1020 1880 -1000
rect 1900 -1020 1920 -1000
rect 1940 -1020 1960 -1000
rect 1980 -1020 2000 -1000
rect 2020 -1020 2040 -1000
rect 2060 -1020 2080 -1000
rect 2100 -1020 2120 -1000
rect 2140 -1020 2160 -1000
rect 2180 -1020 2200 -1000
rect 2220 -1020 2240 -1000
rect 2260 -1020 2280 -1000
rect 2300 -1020 2320 -1000
rect 2340 -1020 2360 -1000
rect 2380 -1020 2400 -1000
rect 2420 -1020 2440 -1000
rect 2460 -1020 2480 -1000
rect 2500 -1020 2520 -1000
rect 2540 -1020 2560 -1000
rect 2590 -1020 2605 -1000
rect 105 -1030 2605 -1020
rect -70 -1045 85 -1035
rect -70 -1070 -60 -1045
rect -40 -1070 -20 -1045
rect 0 -1070 20 -1045
rect 40 -1070 60 -1045
rect -70 -1080 85 -1070
rect 105 -1095 2605 -1085
rect 105 -1115 120 -1095
rect 140 -1115 160 -1095
rect 180 -1115 200 -1095
rect 220 -1115 240 -1095
rect 260 -1115 280 -1095
rect 300 -1115 320 -1095
rect 340 -1115 360 -1095
rect 380 -1115 400 -1095
rect 420 -1115 440 -1095
rect 460 -1115 480 -1095
rect 500 -1115 520 -1095
rect 540 -1115 560 -1095
rect 580 -1115 600 -1095
rect 620 -1115 640 -1095
rect 660 -1115 680 -1095
rect 700 -1115 720 -1095
rect 740 -1115 760 -1095
rect 780 -1115 800 -1095
rect 820 -1115 840 -1095
rect 860 -1115 880 -1095
rect 900 -1115 920 -1095
rect 940 -1115 960 -1095
rect 980 -1115 1000 -1095
rect 1020 -1115 1040 -1095
rect 1060 -1115 1080 -1095
rect 1100 -1115 1120 -1095
rect 1140 -1115 1160 -1095
rect 1180 -1115 1200 -1095
rect 1220 -1115 1240 -1095
rect 1260 -1115 1280 -1095
rect 1300 -1115 1320 -1095
rect 1340 -1115 1360 -1095
rect 1380 -1115 1400 -1095
rect 1420 -1115 1440 -1095
rect 1460 -1115 1480 -1095
rect 1500 -1115 1520 -1095
rect 1540 -1115 1560 -1095
rect 1580 -1115 1600 -1095
rect 1620 -1115 1640 -1095
rect 1660 -1115 1680 -1095
rect 1700 -1115 1720 -1095
rect 1740 -1115 1760 -1095
rect 1780 -1115 1800 -1095
rect 1820 -1115 1840 -1095
rect 1860 -1115 1880 -1095
rect 1900 -1115 1920 -1095
rect 1940 -1115 1960 -1095
rect 1980 -1115 2000 -1095
rect 2020 -1115 2040 -1095
rect 2060 -1115 2080 -1095
rect 2100 -1115 2120 -1095
rect 2140 -1115 2160 -1095
rect 2180 -1115 2200 -1095
rect 2220 -1115 2240 -1095
rect 2260 -1115 2280 -1095
rect 2300 -1115 2320 -1095
rect 2340 -1115 2360 -1095
rect 2380 -1115 2400 -1095
rect 2420 -1115 2440 -1095
rect 2460 -1115 2480 -1095
rect 2500 -1115 2520 -1095
rect 2540 -1115 2560 -1095
rect 2590 -1115 2605 -1095
rect 105 -1125 2605 -1115
rect -70 -1140 85 -1130
rect -70 -1165 -60 -1140
rect -40 -1165 -20 -1140
rect 0 -1165 20 -1140
rect 40 -1165 60 -1140
rect -70 -1175 85 -1165
rect 105 -1190 2605 -1180
rect 105 -1210 120 -1190
rect 140 -1210 160 -1190
rect 180 -1210 200 -1190
rect 220 -1210 240 -1190
rect 260 -1210 280 -1190
rect 300 -1210 320 -1190
rect 340 -1210 360 -1190
rect 380 -1210 400 -1190
rect 420 -1210 440 -1190
rect 460 -1210 480 -1190
rect 500 -1210 520 -1190
rect 540 -1210 560 -1190
rect 580 -1210 600 -1190
rect 620 -1210 640 -1190
rect 660 -1210 680 -1190
rect 700 -1210 720 -1190
rect 740 -1210 760 -1190
rect 780 -1210 800 -1190
rect 820 -1210 840 -1190
rect 860 -1210 880 -1190
rect 900 -1210 920 -1190
rect 940 -1210 960 -1190
rect 980 -1210 1000 -1190
rect 1020 -1210 1040 -1190
rect 1060 -1210 1080 -1190
rect 1100 -1210 1120 -1190
rect 1140 -1210 1160 -1190
rect 1180 -1210 1200 -1190
rect 1220 -1210 1240 -1190
rect 1260 -1210 1280 -1190
rect 1300 -1210 1320 -1190
rect 1340 -1210 1360 -1190
rect 1380 -1210 1400 -1190
rect 1420 -1210 1440 -1190
rect 1460 -1210 1480 -1190
rect 1500 -1210 1520 -1190
rect 1540 -1210 1560 -1190
rect 1580 -1210 1600 -1190
rect 1620 -1210 1640 -1190
rect 1660 -1210 1680 -1190
rect 1700 -1210 1720 -1190
rect 1740 -1210 1760 -1190
rect 1780 -1210 1800 -1190
rect 1820 -1210 1840 -1190
rect 1860 -1210 1880 -1190
rect 1900 -1210 1920 -1190
rect 1940 -1210 1960 -1190
rect 1980 -1210 2000 -1190
rect 2020 -1210 2040 -1190
rect 2060 -1210 2080 -1190
rect 2100 -1210 2120 -1190
rect 2140 -1210 2160 -1190
rect 2180 -1210 2200 -1190
rect 2220 -1210 2240 -1190
rect 2260 -1210 2280 -1190
rect 2300 -1210 2320 -1190
rect 2340 -1210 2360 -1190
rect 2380 -1210 2400 -1190
rect 2420 -1210 2440 -1190
rect 2460 -1210 2480 -1190
rect 2500 -1210 2520 -1190
rect 2540 -1210 2560 -1190
rect 2590 -1210 2605 -1190
rect 105 -1220 2605 -1210
rect -70 -1235 85 -1225
rect -70 -1260 -60 -1235
rect -40 -1260 -20 -1235
rect 0 -1260 20 -1235
rect 40 -1260 60 -1235
rect -70 -1270 85 -1260
rect 105 -1285 2605 -1275
rect 105 -1305 120 -1285
rect 140 -1305 160 -1285
rect 180 -1305 200 -1285
rect 220 -1305 240 -1285
rect 260 -1305 280 -1285
rect 300 -1305 320 -1285
rect 340 -1305 360 -1285
rect 380 -1305 400 -1285
rect 420 -1305 440 -1285
rect 460 -1305 480 -1285
rect 500 -1305 520 -1285
rect 540 -1305 560 -1285
rect 580 -1305 600 -1285
rect 620 -1305 640 -1285
rect 660 -1305 680 -1285
rect 700 -1305 720 -1285
rect 740 -1305 760 -1285
rect 780 -1305 800 -1285
rect 820 -1305 840 -1285
rect 860 -1305 880 -1285
rect 900 -1305 920 -1285
rect 940 -1305 960 -1285
rect 980 -1305 1000 -1285
rect 1020 -1305 1040 -1285
rect 1060 -1305 1080 -1285
rect 1100 -1305 1120 -1285
rect 1140 -1305 1160 -1285
rect 1180 -1305 1200 -1285
rect 1220 -1305 1240 -1285
rect 1260 -1305 1280 -1285
rect 1300 -1305 1320 -1285
rect 1340 -1305 1360 -1285
rect 1380 -1305 1400 -1285
rect 1420 -1305 1440 -1285
rect 1460 -1305 1480 -1285
rect 1500 -1305 1520 -1285
rect 1540 -1305 1560 -1285
rect 1580 -1305 1600 -1285
rect 1620 -1305 1640 -1285
rect 1660 -1305 1680 -1285
rect 1700 -1305 1720 -1285
rect 1740 -1305 1760 -1285
rect 1780 -1305 1800 -1285
rect 1820 -1305 1840 -1285
rect 1860 -1305 1880 -1285
rect 1900 -1305 1920 -1285
rect 1940 -1305 1960 -1285
rect 1980 -1305 2000 -1285
rect 2020 -1305 2040 -1285
rect 2060 -1305 2080 -1285
rect 2100 -1305 2120 -1285
rect 2140 -1305 2160 -1285
rect 2180 -1305 2200 -1285
rect 2220 -1305 2240 -1285
rect 2260 -1305 2280 -1285
rect 2300 -1305 2320 -1285
rect 2340 -1305 2360 -1285
rect 2380 -1305 2400 -1285
rect 2420 -1305 2440 -1285
rect 2460 -1305 2480 -1285
rect 2500 -1305 2520 -1285
rect 2540 -1305 2560 -1285
rect 2590 -1305 2605 -1285
rect 105 -1315 2605 -1305
rect -70 -1330 85 -1320
rect -70 -1355 -60 -1330
rect -40 -1355 -20 -1330
rect 0 -1355 20 -1330
rect 40 -1355 60 -1330
rect -70 -1365 85 -1355
rect 105 -1380 2605 -1370
rect 105 -1400 120 -1380
rect 140 -1400 160 -1380
rect 180 -1400 200 -1380
rect 220 -1400 240 -1380
rect 260 -1400 280 -1380
rect 300 -1400 320 -1380
rect 340 -1400 360 -1380
rect 380 -1400 400 -1380
rect 420 -1400 440 -1380
rect 460 -1400 480 -1380
rect 500 -1400 520 -1380
rect 540 -1400 560 -1380
rect 580 -1400 600 -1380
rect 620 -1400 640 -1380
rect 660 -1400 680 -1380
rect 700 -1400 720 -1380
rect 740 -1400 760 -1380
rect 780 -1400 800 -1380
rect 820 -1400 840 -1380
rect 860 -1400 880 -1380
rect 900 -1400 920 -1380
rect 940 -1400 960 -1380
rect 980 -1400 1000 -1380
rect 1020 -1400 1040 -1380
rect 1060 -1400 1080 -1380
rect 1100 -1400 1120 -1380
rect 1140 -1400 1160 -1380
rect 1180 -1400 1200 -1380
rect 1220 -1400 1240 -1380
rect 1260 -1400 1280 -1380
rect 1300 -1400 1320 -1380
rect 1340 -1400 1360 -1380
rect 1380 -1400 1400 -1380
rect 1420 -1400 1440 -1380
rect 1460 -1400 1480 -1380
rect 1500 -1400 1520 -1380
rect 1540 -1400 1560 -1380
rect 1580 -1400 1600 -1380
rect 1620 -1400 1640 -1380
rect 1660 -1400 1680 -1380
rect 1700 -1400 1720 -1380
rect 1740 -1400 1760 -1380
rect 1780 -1400 1800 -1380
rect 1820 -1400 1840 -1380
rect 1860 -1400 1880 -1380
rect 1900 -1400 1920 -1380
rect 1940 -1400 1960 -1380
rect 1980 -1400 2000 -1380
rect 2020 -1400 2040 -1380
rect 2060 -1400 2080 -1380
rect 2100 -1400 2120 -1380
rect 2140 -1400 2160 -1380
rect 2180 -1400 2200 -1380
rect 2220 -1400 2240 -1380
rect 2260 -1400 2280 -1380
rect 2300 -1400 2320 -1380
rect 2340 -1400 2360 -1380
rect 2380 -1400 2400 -1380
rect 2420 -1400 2440 -1380
rect 2460 -1400 2480 -1380
rect 2500 -1400 2520 -1380
rect 2540 -1400 2560 -1380
rect 2590 -1400 2605 -1380
rect 105 -1410 2605 -1400
rect -70 -1425 85 -1415
rect -70 -1450 -60 -1425
rect -40 -1450 -20 -1425
rect 0 -1450 20 -1425
rect 40 -1450 60 -1425
rect -70 -1460 85 -1450
rect 105 -1475 2605 -1465
rect 105 -1495 120 -1475
rect 140 -1495 160 -1475
rect 180 -1495 200 -1475
rect 220 -1495 240 -1475
rect 260 -1495 280 -1475
rect 300 -1495 320 -1475
rect 340 -1495 360 -1475
rect 380 -1495 400 -1475
rect 420 -1495 440 -1475
rect 460 -1495 480 -1475
rect 500 -1495 520 -1475
rect 540 -1495 560 -1475
rect 580 -1495 600 -1475
rect 620 -1495 640 -1475
rect 660 -1495 680 -1475
rect 700 -1495 720 -1475
rect 740 -1495 760 -1475
rect 780 -1495 800 -1475
rect 820 -1495 840 -1475
rect 860 -1495 880 -1475
rect 900 -1495 920 -1475
rect 940 -1495 960 -1475
rect 980 -1495 1000 -1475
rect 1020 -1495 1040 -1475
rect 1060 -1495 1080 -1475
rect 1100 -1495 1120 -1475
rect 1140 -1495 1160 -1475
rect 1180 -1495 1200 -1475
rect 1220 -1495 1240 -1475
rect 1260 -1495 1280 -1475
rect 1300 -1495 1320 -1475
rect 1340 -1495 1360 -1475
rect 1380 -1495 1400 -1475
rect 1420 -1495 1440 -1475
rect 1460 -1495 1480 -1475
rect 1500 -1495 1520 -1475
rect 1540 -1495 1560 -1475
rect 1580 -1495 1600 -1475
rect 1620 -1495 1640 -1475
rect 1660 -1495 1680 -1475
rect 1700 -1495 1720 -1475
rect 1740 -1495 1760 -1475
rect 1780 -1495 1800 -1475
rect 1820 -1495 1840 -1475
rect 1860 -1495 1880 -1475
rect 1900 -1495 1920 -1475
rect 1940 -1495 1960 -1475
rect 1980 -1495 2000 -1475
rect 2020 -1495 2040 -1475
rect 2060 -1495 2080 -1475
rect 2100 -1495 2120 -1475
rect 2140 -1495 2160 -1475
rect 2180 -1495 2200 -1475
rect 2220 -1495 2240 -1475
rect 2260 -1495 2280 -1475
rect 2300 -1495 2320 -1475
rect 2340 -1495 2360 -1475
rect 2380 -1495 2400 -1475
rect 2420 -1495 2440 -1475
rect 2460 -1495 2480 -1475
rect 2500 -1495 2520 -1475
rect 2540 -1495 2560 -1475
rect 2590 -1495 2605 -1475
rect 105 -1505 2605 -1495
rect -70 -1520 85 -1510
rect -70 -1545 -60 -1520
rect -40 -1545 -20 -1520
rect 0 -1545 20 -1520
rect 40 -1545 60 -1520
rect -70 -1555 85 -1545
rect 105 -1570 2605 -1560
rect 105 -1590 120 -1570
rect 140 -1590 160 -1570
rect 180 -1590 200 -1570
rect 220 -1590 240 -1570
rect 260 -1590 280 -1570
rect 300 -1590 320 -1570
rect 340 -1590 360 -1570
rect 380 -1590 400 -1570
rect 420 -1590 440 -1570
rect 460 -1590 480 -1570
rect 500 -1590 520 -1570
rect 540 -1590 560 -1570
rect 580 -1590 600 -1570
rect 620 -1590 640 -1570
rect 660 -1590 680 -1570
rect 700 -1590 720 -1570
rect 740 -1590 760 -1570
rect 780 -1590 800 -1570
rect 820 -1590 840 -1570
rect 860 -1590 880 -1570
rect 900 -1590 920 -1570
rect 940 -1590 960 -1570
rect 980 -1590 1000 -1570
rect 1020 -1590 1040 -1570
rect 1060 -1590 1080 -1570
rect 1100 -1590 1120 -1570
rect 1140 -1590 1160 -1570
rect 1180 -1590 1200 -1570
rect 1220 -1590 1240 -1570
rect 1260 -1590 1280 -1570
rect 1300 -1590 1320 -1570
rect 1340 -1590 1360 -1570
rect 1380 -1590 1400 -1570
rect 1420 -1590 1440 -1570
rect 1460 -1590 1480 -1570
rect 1500 -1590 1520 -1570
rect 1540 -1590 1560 -1570
rect 1580 -1590 1600 -1570
rect 1620 -1590 1640 -1570
rect 1660 -1590 1680 -1570
rect 1700 -1590 1720 -1570
rect 1740 -1590 1760 -1570
rect 1780 -1590 1800 -1570
rect 1820 -1590 1840 -1570
rect 1860 -1590 1880 -1570
rect 1900 -1590 1920 -1570
rect 1940 -1590 1960 -1570
rect 1980 -1590 2000 -1570
rect 2020 -1590 2040 -1570
rect 2060 -1590 2080 -1570
rect 2100 -1590 2120 -1570
rect 2140 -1590 2160 -1570
rect 2180 -1590 2200 -1570
rect 2220 -1590 2240 -1570
rect 2260 -1590 2280 -1570
rect 2300 -1590 2320 -1570
rect 2340 -1590 2360 -1570
rect 2380 -1590 2400 -1570
rect 2420 -1590 2440 -1570
rect 2460 -1590 2480 -1570
rect 2500 -1590 2520 -1570
rect 2540 -1590 2560 -1570
rect 2590 -1590 2605 -1570
rect 105 -1600 2605 -1590
rect -70 -1615 85 -1605
rect -70 -1640 -60 -1615
rect -40 -1640 -20 -1615
rect 0 -1640 20 -1615
rect 40 -1640 60 -1615
rect -70 -1650 85 -1640
rect 105 -1665 2605 -1655
rect 105 -1685 120 -1665
rect 140 -1685 160 -1665
rect 180 -1685 200 -1665
rect 220 -1685 240 -1665
rect 260 -1685 280 -1665
rect 300 -1685 320 -1665
rect 340 -1685 360 -1665
rect 380 -1685 400 -1665
rect 420 -1685 440 -1665
rect 460 -1685 480 -1665
rect 500 -1685 520 -1665
rect 540 -1685 560 -1665
rect 580 -1685 600 -1665
rect 620 -1685 640 -1665
rect 660 -1685 680 -1665
rect 700 -1685 720 -1665
rect 740 -1685 760 -1665
rect 780 -1685 800 -1665
rect 820 -1685 840 -1665
rect 860 -1685 880 -1665
rect 900 -1685 920 -1665
rect 940 -1685 960 -1665
rect 980 -1685 1000 -1665
rect 1020 -1685 1040 -1665
rect 1060 -1685 1080 -1665
rect 1100 -1685 1120 -1665
rect 1140 -1685 1160 -1665
rect 1180 -1685 1200 -1665
rect 1220 -1685 1240 -1665
rect 1260 -1685 1280 -1665
rect 1300 -1685 1320 -1665
rect 1340 -1685 1360 -1665
rect 1380 -1685 1400 -1665
rect 1420 -1685 1440 -1665
rect 1460 -1685 1480 -1665
rect 1500 -1685 1520 -1665
rect 1540 -1685 1560 -1665
rect 1580 -1685 1600 -1665
rect 1620 -1685 1640 -1665
rect 1660 -1685 1680 -1665
rect 1700 -1685 1720 -1665
rect 1740 -1685 1760 -1665
rect 1780 -1685 1800 -1665
rect 1820 -1685 1840 -1665
rect 1860 -1685 1880 -1665
rect 1900 -1685 1920 -1665
rect 1940 -1685 1960 -1665
rect 1980 -1685 2000 -1665
rect 2020 -1685 2040 -1665
rect 2060 -1685 2080 -1665
rect 2100 -1685 2120 -1665
rect 2140 -1685 2160 -1665
rect 2180 -1685 2200 -1665
rect 2220 -1685 2240 -1665
rect 2260 -1685 2280 -1665
rect 2300 -1685 2320 -1665
rect 2340 -1685 2360 -1665
rect 2380 -1685 2400 -1665
rect 2420 -1685 2440 -1665
rect 2460 -1685 2480 -1665
rect 2500 -1685 2520 -1665
rect 2540 -1685 2560 -1665
rect 2590 -1685 2605 -1665
rect 105 -1695 2605 -1685
rect -70 -1710 85 -1700
rect -70 -1735 -60 -1710
rect -40 -1735 -20 -1710
rect 0 -1735 20 -1710
rect 40 -1735 60 -1710
rect -70 -1745 85 -1735
rect 105 -1760 2605 -1750
rect 105 -1780 120 -1760
rect 140 -1780 160 -1760
rect 180 -1780 200 -1760
rect 220 -1780 240 -1760
rect 260 -1780 280 -1760
rect 300 -1780 320 -1760
rect 340 -1780 360 -1760
rect 380 -1780 400 -1760
rect 420 -1780 440 -1760
rect 460 -1780 480 -1760
rect 500 -1780 520 -1760
rect 540 -1780 560 -1760
rect 580 -1780 600 -1760
rect 620 -1780 640 -1760
rect 660 -1780 680 -1760
rect 700 -1780 720 -1760
rect 740 -1780 760 -1760
rect 780 -1780 800 -1760
rect 820 -1780 840 -1760
rect 860 -1780 880 -1760
rect 900 -1780 920 -1760
rect 940 -1780 960 -1760
rect 980 -1780 1000 -1760
rect 1020 -1780 1040 -1760
rect 1060 -1780 1080 -1760
rect 1100 -1780 1120 -1760
rect 1140 -1780 1160 -1760
rect 1180 -1780 1200 -1760
rect 1220 -1780 1240 -1760
rect 1260 -1780 1280 -1760
rect 1300 -1780 1320 -1760
rect 1340 -1780 1360 -1760
rect 1380 -1780 1400 -1760
rect 1420 -1780 1440 -1760
rect 1460 -1780 1480 -1760
rect 1500 -1780 1520 -1760
rect 1540 -1780 1560 -1760
rect 1580 -1780 1600 -1760
rect 1620 -1780 1640 -1760
rect 1660 -1780 1680 -1760
rect 1700 -1780 1720 -1760
rect 1740 -1780 1760 -1760
rect 1780 -1780 1800 -1760
rect 1820 -1780 1840 -1760
rect 1860 -1780 1880 -1760
rect 1900 -1780 1920 -1760
rect 1940 -1780 1960 -1760
rect 1980 -1780 2000 -1760
rect 2020 -1780 2040 -1760
rect 2060 -1780 2080 -1760
rect 2100 -1780 2120 -1760
rect 2140 -1780 2160 -1760
rect 2180 -1780 2200 -1760
rect 2220 -1780 2240 -1760
rect 2260 -1780 2280 -1760
rect 2300 -1780 2320 -1760
rect 2340 -1780 2360 -1760
rect 2380 -1780 2400 -1760
rect 2420 -1780 2440 -1760
rect 2460 -1780 2480 -1760
rect 2500 -1780 2520 -1760
rect 2540 -1780 2560 -1760
rect 2590 -1780 2605 -1760
rect 105 -1790 2605 -1780
rect -70 -1805 85 -1795
rect -70 -1830 -60 -1805
rect -40 -1830 -20 -1805
rect 0 -1830 20 -1805
rect 40 -1830 60 -1805
rect -70 -1840 85 -1830
rect 105 -1855 2605 -1845
rect 105 -1875 120 -1855
rect 140 -1875 160 -1855
rect 180 -1875 200 -1855
rect 220 -1875 240 -1855
rect 260 -1875 280 -1855
rect 300 -1875 320 -1855
rect 340 -1875 360 -1855
rect 380 -1875 400 -1855
rect 420 -1875 440 -1855
rect 460 -1875 480 -1855
rect 500 -1875 520 -1855
rect 540 -1875 560 -1855
rect 580 -1875 600 -1855
rect 620 -1875 640 -1855
rect 660 -1875 680 -1855
rect 700 -1875 720 -1855
rect 740 -1875 760 -1855
rect 780 -1875 800 -1855
rect 820 -1875 840 -1855
rect 860 -1875 880 -1855
rect 900 -1875 920 -1855
rect 940 -1875 960 -1855
rect 980 -1875 1000 -1855
rect 1020 -1875 1040 -1855
rect 1060 -1875 1080 -1855
rect 1100 -1875 1120 -1855
rect 1140 -1875 1160 -1855
rect 1180 -1875 1200 -1855
rect 1220 -1875 1240 -1855
rect 1260 -1875 1280 -1855
rect 1300 -1875 1320 -1855
rect 1340 -1875 1360 -1855
rect 1380 -1875 1400 -1855
rect 1420 -1875 1440 -1855
rect 1460 -1875 1480 -1855
rect 1500 -1875 1520 -1855
rect 1540 -1875 1560 -1855
rect 1580 -1875 1600 -1855
rect 1620 -1875 1640 -1855
rect 1660 -1875 1680 -1855
rect 1700 -1875 1720 -1855
rect 1740 -1875 1760 -1855
rect 1780 -1875 1800 -1855
rect 1820 -1875 1840 -1855
rect 1860 -1875 1880 -1855
rect 1900 -1875 1920 -1855
rect 1940 -1875 1960 -1855
rect 1980 -1875 2000 -1855
rect 2020 -1875 2040 -1855
rect 2060 -1875 2080 -1855
rect 2100 -1875 2120 -1855
rect 2140 -1875 2160 -1855
rect 2180 -1875 2200 -1855
rect 2220 -1875 2240 -1855
rect 2260 -1875 2280 -1855
rect 2300 -1875 2320 -1855
rect 2340 -1875 2360 -1855
rect 2380 -1875 2400 -1855
rect 2420 -1875 2440 -1855
rect 2460 -1875 2480 -1855
rect 2500 -1875 2520 -1855
rect 2540 -1875 2560 -1855
rect 2590 -1875 2605 -1855
rect 105 -1885 2605 -1875
rect -70 -1900 85 -1890
rect -70 -1925 -60 -1900
rect -40 -1925 -20 -1900
rect 0 -1925 20 -1900
rect 40 -1925 60 -1900
rect -70 -1935 85 -1925
rect 105 -1950 2605 -1940
rect 105 -1970 120 -1950
rect 140 -1970 160 -1950
rect 180 -1970 200 -1950
rect 220 -1970 240 -1950
rect 260 -1970 280 -1950
rect 300 -1970 320 -1950
rect 340 -1970 360 -1950
rect 380 -1970 400 -1950
rect 420 -1970 440 -1950
rect 460 -1970 480 -1950
rect 500 -1970 520 -1950
rect 540 -1970 560 -1950
rect 580 -1970 600 -1950
rect 620 -1970 640 -1950
rect 660 -1970 680 -1950
rect 700 -1970 720 -1950
rect 740 -1970 760 -1950
rect 780 -1970 800 -1950
rect 820 -1970 840 -1950
rect 860 -1970 880 -1950
rect 900 -1970 920 -1950
rect 940 -1970 960 -1950
rect 980 -1970 1000 -1950
rect 1020 -1970 1040 -1950
rect 1060 -1970 1080 -1950
rect 1100 -1970 1120 -1950
rect 1140 -1970 1160 -1950
rect 1180 -1970 1200 -1950
rect 1220 -1970 1240 -1950
rect 1260 -1970 1280 -1950
rect 1300 -1970 1320 -1950
rect 1340 -1970 1360 -1950
rect 1380 -1970 1400 -1950
rect 1420 -1970 1440 -1950
rect 1460 -1970 1480 -1950
rect 1500 -1970 1520 -1950
rect 1540 -1970 1560 -1950
rect 1580 -1970 1600 -1950
rect 1620 -1970 1640 -1950
rect 1660 -1970 1680 -1950
rect 1700 -1970 1720 -1950
rect 1740 -1970 1760 -1950
rect 1780 -1970 1800 -1950
rect 1820 -1970 1840 -1950
rect 1860 -1970 1880 -1950
rect 1900 -1970 1920 -1950
rect 1940 -1970 1960 -1950
rect 1980 -1970 2000 -1950
rect 2020 -1970 2040 -1950
rect 2060 -1970 2080 -1950
rect 2100 -1970 2120 -1950
rect 2140 -1970 2160 -1950
rect 2180 -1970 2200 -1950
rect 2220 -1970 2240 -1950
rect 2260 -1970 2280 -1950
rect 2300 -1970 2320 -1950
rect 2340 -1970 2360 -1950
rect 2380 -1970 2400 -1950
rect 2420 -1970 2440 -1950
rect 2460 -1970 2480 -1950
rect 2500 -1970 2520 -1950
rect 2540 -1970 2560 -1950
rect 2590 -1970 2605 -1950
rect 105 -1980 2605 -1970
rect -70 -1995 85 -1985
rect -70 -2020 -60 -1995
rect -40 -2020 -20 -1995
rect 0 -2020 20 -1995
rect 40 -2020 60 -1995
rect -70 -2030 85 -2020
rect 105 -2045 2605 -2035
rect 105 -2065 120 -2045
rect 140 -2065 160 -2045
rect 180 -2065 200 -2045
rect 220 -2065 240 -2045
rect 260 -2065 280 -2045
rect 300 -2065 320 -2045
rect 340 -2065 360 -2045
rect 380 -2065 400 -2045
rect 420 -2065 440 -2045
rect 460 -2065 480 -2045
rect 500 -2065 520 -2045
rect 540 -2065 560 -2045
rect 580 -2065 600 -2045
rect 620 -2065 640 -2045
rect 660 -2065 680 -2045
rect 700 -2065 720 -2045
rect 740 -2065 760 -2045
rect 780 -2065 800 -2045
rect 820 -2065 840 -2045
rect 860 -2065 880 -2045
rect 900 -2065 920 -2045
rect 940 -2065 960 -2045
rect 980 -2065 1000 -2045
rect 1020 -2065 1040 -2045
rect 1060 -2065 1080 -2045
rect 1100 -2065 1120 -2045
rect 1140 -2065 1160 -2045
rect 1180 -2065 1200 -2045
rect 1220 -2065 1240 -2045
rect 1260 -2065 1280 -2045
rect 1300 -2065 1320 -2045
rect 1340 -2065 1360 -2045
rect 1380 -2065 1400 -2045
rect 1420 -2065 1440 -2045
rect 1460 -2065 1480 -2045
rect 1500 -2065 1520 -2045
rect 1540 -2065 1560 -2045
rect 1580 -2065 1600 -2045
rect 1620 -2065 1640 -2045
rect 1660 -2065 1680 -2045
rect 1700 -2065 1720 -2045
rect 1740 -2065 1760 -2045
rect 1780 -2065 1800 -2045
rect 1820 -2065 1840 -2045
rect 1860 -2065 1880 -2045
rect 1900 -2065 1920 -2045
rect 1940 -2065 1960 -2045
rect 1980 -2065 2000 -2045
rect 2020 -2065 2040 -2045
rect 2060 -2065 2080 -2045
rect 2100 -2065 2120 -2045
rect 2140 -2065 2160 -2045
rect 2180 -2065 2200 -2045
rect 2220 -2065 2240 -2045
rect 2260 -2065 2280 -2045
rect 2300 -2065 2320 -2045
rect 2340 -2065 2360 -2045
rect 2380 -2065 2400 -2045
rect 2420 -2065 2440 -2045
rect 2460 -2065 2480 -2045
rect 2500 -2065 2520 -2045
rect 2540 -2065 2560 -2045
rect 2590 -2065 2605 -2045
rect 105 -2075 2605 -2065
rect -70 -2090 85 -2080
rect -70 -2115 -60 -2090
rect -40 -2115 -20 -2090
rect 0 -2115 20 -2090
rect 40 -2115 60 -2090
rect -70 -2125 85 -2115
rect 105 -2140 2605 -2130
rect 105 -2160 120 -2140
rect 140 -2160 160 -2140
rect 180 -2160 200 -2140
rect 220 -2160 240 -2140
rect 260 -2160 280 -2140
rect 300 -2160 320 -2140
rect 340 -2160 360 -2140
rect 380 -2160 400 -2140
rect 420 -2160 440 -2140
rect 460 -2160 480 -2140
rect 500 -2160 520 -2140
rect 540 -2160 560 -2140
rect 580 -2160 600 -2140
rect 620 -2160 640 -2140
rect 660 -2160 680 -2140
rect 700 -2160 720 -2140
rect 740 -2160 760 -2140
rect 780 -2160 800 -2140
rect 820 -2160 840 -2140
rect 860 -2160 880 -2140
rect 900 -2160 920 -2140
rect 940 -2160 960 -2140
rect 980 -2160 1000 -2140
rect 1020 -2160 1040 -2140
rect 1060 -2160 1080 -2140
rect 1100 -2160 1120 -2140
rect 1140 -2160 1160 -2140
rect 1180 -2160 1200 -2140
rect 1220 -2160 1240 -2140
rect 1260 -2160 1280 -2140
rect 1300 -2160 1320 -2140
rect 1340 -2160 1360 -2140
rect 1380 -2160 1400 -2140
rect 1420 -2160 1440 -2140
rect 1460 -2160 1480 -2140
rect 1500 -2160 1520 -2140
rect 1540 -2160 1560 -2140
rect 1580 -2160 1600 -2140
rect 1620 -2160 1640 -2140
rect 1660 -2160 1680 -2140
rect 1700 -2160 1720 -2140
rect 1740 -2160 1760 -2140
rect 1780 -2160 1800 -2140
rect 1820 -2160 1840 -2140
rect 1860 -2160 1880 -2140
rect 1900 -2160 1920 -2140
rect 1940 -2160 1960 -2140
rect 1980 -2160 2000 -2140
rect 2020 -2160 2040 -2140
rect 2060 -2160 2080 -2140
rect 2100 -2160 2120 -2140
rect 2140 -2160 2160 -2140
rect 2180 -2160 2200 -2140
rect 2220 -2160 2240 -2140
rect 2260 -2160 2280 -2140
rect 2300 -2160 2320 -2140
rect 2340 -2160 2360 -2140
rect 2380 -2160 2400 -2140
rect 2420 -2160 2440 -2140
rect 2460 -2160 2480 -2140
rect 2500 -2160 2520 -2140
rect 2540 -2160 2560 -2140
rect 2590 -2160 2605 -2140
rect 105 -2170 2605 -2160
rect -70 -2185 85 -2175
rect -70 -2210 -60 -2185
rect -40 -2210 -20 -2185
rect 0 -2210 20 -2185
rect 40 -2210 60 -2185
rect -70 -2220 85 -2210
rect 105 -2235 2605 -2225
rect 105 -2255 120 -2235
rect 140 -2255 160 -2235
rect 180 -2255 200 -2235
rect 220 -2255 240 -2235
rect 260 -2255 280 -2235
rect 300 -2255 320 -2235
rect 340 -2255 360 -2235
rect 380 -2255 400 -2235
rect 420 -2255 440 -2235
rect 460 -2255 480 -2235
rect 500 -2255 520 -2235
rect 540 -2255 560 -2235
rect 580 -2255 600 -2235
rect 620 -2255 640 -2235
rect 660 -2255 680 -2235
rect 700 -2255 720 -2235
rect 740 -2255 760 -2235
rect 780 -2255 800 -2235
rect 820 -2255 840 -2235
rect 860 -2255 880 -2235
rect 900 -2255 920 -2235
rect 940 -2255 960 -2235
rect 980 -2255 1000 -2235
rect 1020 -2255 1040 -2235
rect 1060 -2255 1080 -2235
rect 1100 -2255 1120 -2235
rect 1140 -2255 1160 -2235
rect 1180 -2255 1200 -2235
rect 1220 -2255 1240 -2235
rect 1260 -2255 1280 -2235
rect 1300 -2255 1320 -2235
rect 1340 -2255 1360 -2235
rect 1380 -2255 1400 -2235
rect 1420 -2255 1440 -2235
rect 1460 -2255 1480 -2235
rect 1500 -2255 1520 -2235
rect 1540 -2255 1560 -2235
rect 1580 -2255 1600 -2235
rect 1620 -2255 1640 -2235
rect 1660 -2255 1680 -2235
rect 1700 -2255 1720 -2235
rect 1740 -2255 1760 -2235
rect 1780 -2255 1800 -2235
rect 1820 -2255 1840 -2235
rect 1860 -2255 1880 -2235
rect 1900 -2255 1920 -2235
rect 1940 -2255 1960 -2235
rect 1980 -2255 2000 -2235
rect 2020 -2255 2040 -2235
rect 2060 -2255 2080 -2235
rect 2100 -2255 2120 -2235
rect 2140 -2255 2160 -2235
rect 2180 -2255 2200 -2235
rect 2220 -2255 2240 -2235
rect 2260 -2255 2280 -2235
rect 2300 -2255 2320 -2235
rect 2340 -2255 2360 -2235
rect 2380 -2255 2400 -2235
rect 2420 -2255 2440 -2235
rect 2460 -2255 2480 -2235
rect 2500 -2255 2520 -2235
rect 2540 -2255 2560 -2235
rect 2590 -2255 2605 -2235
rect 105 -2265 2605 -2255
rect -70 -2280 85 -2270
rect -70 -2305 -60 -2280
rect -40 -2305 -20 -2280
rect 0 -2305 20 -2280
rect 40 -2305 60 -2280
rect -70 -2315 85 -2305
rect 105 -2330 2605 -2320
rect 105 -2350 120 -2330
rect 140 -2350 160 -2330
rect 180 -2350 200 -2330
rect 220 -2350 240 -2330
rect 260 -2350 280 -2330
rect 300 -2350 320 -2330
rect 340 -2350 360 -2330
rect 380 -2350 400 -2330
rect 420 -2350 440 -2330
rect 460 -2350 480 -2330
rect 500 -2350 520 -2330
rect 540 -2350 560 -2330
rect 580 -2350 600 -2330
rect 620 -2350 640 -2330
rect 660 -2350 680 -2330
rect 700 -2350 720 -2330
rect 740 -2350 760 -2330
rect 780 -2350 800 -2330
rect 820 -2350 840 -2330
rect 860 -2350 880 -2330
rect 900 -2350 920 -2330
rect 940 -2350 960 -2330
rect 980 -2350 1000 -2330
rect 1020 -2350 1040 -2330
rect 1060 -2350 1080 -2330
rect 1100 -2350 1120 -2330
rect 1140 -2350 1160 -2330
rect 1180 -2350 1200 -2330
rect 1220 -2350 1240 -2330
rect 1260 -2350 1280 -2330
rect 1300 -2350 1320 -2330
rect 1340 -2350 1360 -2330
rect 1380 -2350 1400 -2330
rect 1420 -2350 1440 -2330
rect 1460 -2350 1480 -2330
rect 1500 -2350 1520 -2330
rect 1540 -2350 1560 -2330
rect 1580 -2350 1600 -2330
rect 1620 -2350 1640 -2330
rect 1660 -2350 1680 -2330
rect 1700 -2350 1720 -2330
rect 1740 -2350 1760 -2330
rect 1780 -2350 1800 -2330
rect 1820 -2350 1840 -2330
rect 1860 -2350 1880 -2330
rect 1900 -2350 1920 -2330
rect 1940 -2350 1960 -2330
rect 1980 -2350 2000 -2330
rect 2020 -2350 2040 -2330
rect 2060 -2350 2080 -2330
rect 2100 -2350 2120 -2330
rect 2140 -2350 2160 -2330
rect 2180 -2350 2200 -2330
rect 2220 -2350 2240 -2330
rect 2260 -2350 2280 -2330
rect 2300 -2350 2320 -2330
rect 2340 -2350 2360 -2330
rect 2380 -2350 2400 -2330
rect 2420 -2350 2440 -2330
rect 2460 -2350 2480 -2330
rect 2500 -2350 2520 -2330
rect 2540 -2350 2560 -2330
rect 2590 -2350 2605 -2330
rect 105 -2360 2605 -2350
rect -70 -2375 85 -2365
rect -70 -2400 -60 -2375
rect -40 -2400 -20 -2375
rect 0 -2400 20 -2375
rect 40 -2400 60 -2375
rect -70 -2410 85 -2400
rect 105 -2425 2605 -2415
rect 105 -2445 120 -2425
rect 140 -2445 160 -2425
rect 180 -2445 200 -2425
rect 220 -2445 240 -2425
rect 260 -2445 280 -2425
rect 300 -2445 320 -2425
rect 340 -2445 360 -2425
rect 380 -2445 400 -2425
rect 420 -2445 440 -2425
rect 460 -2445 480 -2425
rect 500 -2445 520 -2425
rect 540 -2445 560 -2425
rect 580 -2445 600 -2425
rect 620 -2445 640 -2425
rect 660 -2445 680 -2425
rect 700 -2445 720 -2425
rect 740 -2445 760 -2425
rect 780 -2445 800 -2425
rect 820 -2445 840 -2425
rect 860 -2445 880 -2425
rect 900 -2445 920 -2425
rect 940 -2445 960 -2425
rect 980 -2445 1000 -2425
rect 1020 -2445 1040 -2425
rect 1060 -2445 1080 -2425
rect 1100 -2445 1120 -2425
rect 1140 -2445 1160 -2425
rect 1180 -2445 1200 -2425
rect 1220 -2445 1240 -2425
rect 1260 -2445 1280 -2425
rect 1300 -2445 1320 -2425
rect 1340 -2445 1360 -2425
rect 1380 -2445 1400 -2425
rect 1420 -2445 1440 -2425
rect 1460 -2445 1480 -2425
rect 1500 -2445 1520 -2425
rect 1540 -2445 1560 -2425
rect 1580 -2445 1600 -2425
rect 1620 -2445 1640 -2425
rect 1660 -2445 1680 -2425
rect 1700 -2445 1720 -2425
rect 1740 -2445 1760 -2425
rect 1780 -2445 1800 -2425
rect 1820 -2445 1840 -2425
rect 1860 -2445 1880 -2425
rect 1900 -2445 1920 -2425
rect 1940 -2445 1960 -2425
rect 1980 -2445 2000 -2425
rect 2020 -2445 2040 -2425
rect 2060 -2445 2080 -2425
rect 2100 -2445 2120 -2425
rect 2140 -2445 2160 -2425
rect 2180 -2445 2200 -2425
rect 2220 -2445 2240 -2425
rect 2260 -2445 2280 -2425
rect 2300 -2445 2320 -2425
rect 2340 -2445 2360 -2425
rect 2380 -2445 2400 -2425
rect 2420 -2445 2440 -2425
rect 2460 -2445 2480 -2425
rect 2500 -2445 2520 -2425
rect 2540 -2445 2560 -2425
rect 2590 -2445 2605 -2425
rect 105 -2455 2605 -2445
rect -70 -2470 85 -2460
rect -70 -2495 -60 -2470
rect -40 -2495 -20 -2470
rect 0 -2495 20 -2470
rect 40 -2495 60 -2470
rect -70 -2505 85 -2495
rect 105 -2520 2605 -2510
rect 105 -2540 120 -2520
rect 140 -2540 160 -2520
rect 180 -2540 200 -2520
rect 220 -2540 240 -2520
rect 260 -2540 280 -2520
rect 300 -2540 320 -2520
rect 340 -2540 360 -2520
rect 380 -2540 400 -2520
rect 420 -2540 440 -2520
rect 460 -2540 480 -2520
rect 500 -2540 520 -2520
rect 540 -2540 560 -2520
rect 580 -2540 600 -2520
rect 620 -2540 640 -2520
rect 660 -2540 680 -2520
rect 700 -2540 720 -2520
rect 740 -2540 760 -2520
rect 780 -2540 800 -2520
rect 820 -2540 840 -2520
rect 860 -2540 880 -2520
rect 900 -2540 920 -2520
rect 940 -2540 960 -2520
rect 980 -2540 1000 -2520
rect 1020 -2540 1040 -2520
rect 1060 -2540 1080 -2520
rect 1100 -2540 1120 -2520
rect 1140 -2540 1160 -2520
rect 1180 -2540 1200 -2520
rect 1220 -2540 1240 -2520
rect 1260 -2540 1280 -2520
rect 1300 -2540 1320 -2520
rect 1340 -2540 1360 -2520
rect 1380 -2540 1400 -2520
rect 1420 -2540 1440 -2520
rect 1460 -2540 1480 -2520
rect 1500 -2540 1520 -2520
rect 1540 -2540 1560 -2520
rect 1580 -2540 1600 -2520
rect 1620 -2540 1640 -2520
rect 1660 -2540 1680 -2520
rect 1700 -2540 1720 -2520
rect 1740 -2540 1760 -2520
rect 1780 -2540 1800 -2520
rect 1820 -2540 1840 -2520
rect 1860 -2540 1880 -2520
rect 1900 -2540 1920 -2520
rect 1940 -2540 1960 -2520
rect 1980 -2540 2000 -2520
rect 2020 -2540 2040 -2520
rect 2060 -2540 2080 -2520
rect 2100 -2540 2120 -2520
rect 2140 -2540 2160 -2520
rect 2180 -2540 2200 -2520
rect 2220 -2540 2240 -2520
rect 2260 -2540 2280 -2520
rect 2300 -2540 2320 -2520
rect 2340 -2540 2360 -2520
rect 2380 -2540 2400 -2520
rect 2420 -2540 2440 -2520
rect 2460 -2540 2480 -2520
rect 2500 -2540 2520 -2520
rect 2540 -2540 2560 -2520
rect 2590 -2540 2605 -2520
rect 105 -2560 2605 -2540
rect 105 -2580 120 -2560
rect 140 -2580 160 -2560
rect 180 -2580 200 -2560
rect 220 -2580 240 -2560
rect 260 -2580 280 -2560
rect 300 -2580 320 -2560
rect 340 -2580 360 -2560
rect 380 -2580 400 -2560
rect 420 -2580 440 -2560
rect 460 -2580 480 -2560
rect 500 -2580 520 -2560
rect 540 -2580 560 -2560
rect 580 -2580 600 -2560
rect 620 -2580 640 -2560
rect 660 -2580 680 -2560
rect 700 -2580 720 -2560
rect 740 -2580 760 -2560
rect 780 -2580 800 -2560
rect 820 -2580 840 -2560
rect 860 -2580 880 -2560
rect 900 -2580 920 -2560
rect 940 -2580 960 -2560
rect 980 -2580 1000 -2560
rect 1020 -2580 1040 -2560
rect 1060 -2580 1080 -2560
rect 1100 -2580 1120 -2560
rect 1140 -2580 1160 -2560
rect 1180 -2580 1200 -2560
rect 1220 -2580 1240 -2560
rect 1260 -2580 1280 -2560
rect 1300 -2580 1320 -2560
rect 1340 -2580 1360 -2560
rect 1380 -2580 1400 -2560
rect 1420 -2580 1440 -2560
rect 1460 -2580 1480 -2560
rect 1500 -2580 1520 -2560
rect 1540 -2580 1560 -2560
rect 1580 -2580 1600 -2560
rect 1620 -2580 1640 -2560
rect 1660 -2580 1680 -2560
rect 1700 -2580 1720 -2560
rect 1740 -2580 1760 -2560
rect 1780 -2580 1800 -2560
rect 1820 -2580 1840 -2560
rect 1860 -2580 1880 -2560
rect 1900 -2580 1920 -2560
rect 1940 -2580 1960 -2560
rect 1980 -2580 2000 -2560
rect 2020 -2580 2040 -2560
rect 2060 -2580 2080 -2560
rect 2100 -2580 2120 -2560
rect 2140 -2580 2160 -2560
rect 2180 -2580 2200 -2560
rect 2220 -2580 2240 -2560
rect 2260 -2580 2280 -2560
rect 2300 -2580 2320 -2560
rect 2340 -2580 2360 -2560
rect 2380 -2580 2400 -2560
rect 2420 -2580 2440 -2560
rect 2460 -2580 2480 -2560
rect 2500 -2580 2520 -2560
rect 2540 -2580 2560 -2560
rect 2590 -2580 2605 -2560
rect 105 -2590 2605 -2580
<< viali >>
rect 200 2345 220 2365
rect 240 2345 260 2365
rect 280 2345 300 2365
rect 320 2345 340 2365
rect 360 2345 380 2365
rect 400 2345 420 2365
rect 440 2345 460 2365
rect 480 2345 500 2365
rect 520 2345 540 2365
rect 560 2345 580 2365
rect 600 2345 620 2365
rect 640 2345 660 2365
rect 680 2345 700 2365
rect 720 2345 740 2365
rect 760 2345 780 2365
rect 800 2345 820 2365
rect 840 2345 860 2365
rect 880 2345 900 2365
rect 920 2345 940 2365
rect 960 2345 980 2365
rect 1000 2345 1020 2365
rect 1040 2345 1060 2365
rect 680 2277 700 2297
rect 720 2277 740 2297
rect 760 2277 780 2297
rect 800 2277 820 2297
rect 840 2277 860 2297
rect 880 2277 900 2297
rect 920 2277 940 2297
rect 960 2277 980 2297
rect 1000 2277 1020 2297
rect 1040 2277 1060 2297
rect 1080 2277 1100 2297
rect 1120 2277 1140 2297
rect 1160 2277 1180 2297
rect 1200 2277 1220 2297
rect 1240 2277 1260 2297
rect 1280 2277 1300 2297
rect 1320 2277 1340 2297
rect 1360 2277 1380 2297
rect 1400 2277 1420 2297
rect 1440 2277 1460 2297
rect 10 2235 30 2255
rect 50 2235 70 2255
rect 90 2235 110 2255
rect 130 2235 150 2255
rect 1760 2195 1780 2215
rect 1800 2195 1820 2215
rect 1840 2195 1860 2215
rect 1880 2195 1900 2215
rect 1920 2195 1940 2215
rect 1960 2195 1980 2215
rect 2000 2195 2020 2215
rect 2040 2195 2060 2215
rect 2080 2195 2100 2215
rect 2120 2195 2140 2215
rect 2160 2195 2180 2215
rect 2200 2195 2220 2215
rect 2240 2195 2260 2215
rect 2280 2195 2300 2215
rect 2320 2195 2340 2215
rect 2360 2195 2380 2215
rect 2400 2195 2420 2215
rect 2440 2195 2460 2215
rect 2480 2195 2500 2215
rect 2520 2195 2540 2215
rect 10 2155 30 2175
rect 50 2155 70 2175
rect 90 2155 110 2175
rect 130 2155 150 2175
rect 680 2113 700 2133
rect 720 2113 740 2133
rect 760 2113 780 2133
rect 800 2113 820 2133
rect 840 2113 860 2133
rect 880 2113 900 2133
rect 920 2113 940 2133
rect 960 2113 980 2133
rect 1000 2113 1020 2133
rect 1040 2113 1060 2133
rect 1080 2113 1100 2133
rect 1120 2113 1140 2133
rect 1160 2113 1180 2133
rect 1200 2113 1220 2133
rect 1240 2113 1260 2133
rect 1280 2113 1300 2133
rect 1320 2113 1340 2133
rect 1360 2113 1380 2133
rect 1400 2113 1420 2133
rect 1440 2113 1460 2133
rect 10 2070 30 2090
rect 50 2070 70 2090
rect 90 2070 110 2090
rect 130 2070 150 2090
rect 1760 2031 1780 2051
rect 1800 2031 1820 2051
rect 1840 2031 1860 2051
rect 1880 2031 1900 2051
rect 1920 2031 1940 2051
rect 1960 2031 1980 2051
rect 2000 2031 2020 2051
rect 2040 2031 2060 2051
rect 2080 2031 2100 2051
rect 2120 2031 2140 2051
rect 2160 2031 2180 2051
rect 2200 2031 2220 2051
rect 2240 2031 2260 2051
rect 2280 2031 2300 2051
rect 2320 2031 2340 2051
rect 2360 2031 2380 2051
rect 2400 2031 2420 2051
rect 2440 2031 2460 2051
rect 2480 2031 2500 2051
rect 2520 2031 2540 2051
rect 10 1990 30 2010
rect 50 1990 70 2010
rect 90 1990 110 2010
rect 130 1990 150 2010
rect 680 1949 700 1969
rect 720 1949 740 1969
rect 760 1949 780 1969
rect 800 1949 820 1969
rect 840 1949 860 1969
rect 880 1949 900 1969
rect 920 1949 940 1969
rect 960 1949 980 1969
rect 1000 1949 1020 1969
rect 1040 1949 1060 1969
rect 1080 1949 1100 1969
rect 1120 1949 1140 1969
rect 1160 1949 1180 1969
rect 1200 1949 1220 1969
rect 1240 1949 1260 1969
rect 1280 1949 1300 1969
rect 1320 1949 1340 1969
rect 1360 1949 1380 1969
rect 1400 1949 1420 1969
rect 1440 1949 1460 1969
rect 10 1910 30 1930
rect 50 1910 70 1930
rect 90 1910 110 1930
rect 130 1910 150 1930
rect 1760 1867 1780 1887
rect 1800 1867 1820 1887
rect 1840 1867 1860 1887
rect 1880 1867 1900 1887
rect 1920 1867 1940 1887
rect 1960 1867 1980 1887
rect 2000 1867 2020 1887
rect 2040 1867 2060 1887
rect 2080 1867 2100 1887
rect 2120 1867 2140 1887
rect 2160 1867 2180 1887
rect 2200 1867 2220 1887
rect 2240 1867 2260 1887
rect 2280 1867 2300 1887
rect 2320 1867 2340 1887
rect 2360 1867 2380 1887
rect 2400 1867 2420 1887
rect 2440 1867 2460 1887
rect 2480 1867 2500 1887
rect 2520 1867 2540 1887
rect 10 1825 30 1845
rect 50 1825 70 1845
rect 90 1825 110 1845
rect 130 1825 150 1845
rect 680 1785 700 1805
rect 720 1785 740 1805
rect 760 1785 780 1805
rect 800 1785 820 1805
rect 840 1785 860 1805
rect 880 1785 900 1805
rect 920 1785 940 1805
rect 960 1785 980 1805
rect 1000 1785 1020 1805
rect 1040 1785 1060 1805
rect 1080 1785 1100 1805
rect 1120 1785 1140 1805
rect 1160 1785 1180 1805
rect 1200 1785 1220 1805
rect 1240 1785 1260 1805
rect 1280 1785 1300 1805
rect 1320 1785 1340 1805
rect 1360 1785 1380 1805
rect 1400 1785 1420 1805
rect 1440 1785 1460 1805
rect 10 1745 30 1765
rect 50 1745 70 1765
rect 90 1745 110 1765
rect 130 1745 150 1765
rect 1760 1703 1780 1723
rect 1800 1703 1820 1723
rect 1840 1703 1860 1723
rect 1880 1703 1900 1723
rect 1920 1703 1940 1723
rect 1960 1703 1980 1723
rect 2000 1703 2020 1723
rect 2040 1703 2060 1723
rect 2080 1703 2100 1723
rect 2120 1703 2140 1723
rect 2160 1703 2180 1723
rect 2200 1703 2220 1723
rect 2240 1703 2260 1723
rect 2280 1703 2300 1723
rect 2320 1703 2340 1723
rect 2360 1703 2380 1723
rect 2400 1703 2420 1723
rect 2440 1703 2460 1723
rect 2480 1703 2500 1723
rect 2520 1703 2540 1723
rect 10 1660 30 1680
rect 50 1660 70 1680
rect 90 1660 110 1680
rect 130 1660 150 1680
rect 680 1621 700 1641
rect 720 1621 740 1641
rect 760 1621 780 1641
rect 800 1621 820 1641
rect 840 1621 860 1641
rect 880 1621 900 1641
rect 920 1621 940 1641
rect 960 1621 980 1641
rect 1000 1621 1020 1641
rect 1040 1621 1060 1641
rect 1080 1621 1100 1641
rect 1120 1621 1140 1641
rect 1160 1621 1180 1641
rect 1200 1621 1220 1641
rect 1240 1621 1260 1641
rect 1280 1621 1300 1641
rect 1320 1621 1340 1641
rect 1360 1621 1380 1641
rect 1400 1621 1420 1641
rect 1440 1621 1460 1641
rect 10 1580 30 1600
rect 50 1580 70 1600
rect 90 1580 110 1600
rect 130 1580 150 1600
rect 1760 1539 1780 1559
rect 1800 1539 1820 1559
rect 1840 1539 1860 1559
rect 1880 1539 1900 1559
rect 1920 1539 1940 1559
rect 1960 1539 1980 1559
rect 2000 1539 2020 1559
rect 2040 1539 2060 1559
rect 2080 1539 2100 1559
rect 2120 1539 2140 1559
rect 2160 1539 2180 1559
rect 2200 1539 2220 1559
rect 2240 1539 2260 1559
rect 2280 1539 2300 1559
rect 2320 1539 2340 1559
rect 2360 1539 2380 1559
rect 2400 1539 2420 1559
rect 2440 1539 2460 1559
rect 2480 1539 2500 1559
rect 2520 1539 2540 1559
rect 10 1500 30 1520
rect 50 1500 70 1520
rect 90 1500 110 1520
rect 130 1500 150 1520
rect 680 1457 700 1477
rect 720 1457 740 1477
rect 760 1457 780 1477
rect 800 1457 820 1477
rect 840 1457 860 1477
rect 880 1457 900 1477
rect 920 1457 940 1477
rect 960 1457 980 1477
rect 1000 1457 1020 1477
rect 1040 1457 1060 1477
rect 1080 1457 1100 1477
rect 1120 1457 1140 1477
rect 1160 1457 1180 1477
rect 1200 1457 1220 1477
rect 1240 1457 1260 1477
rect 1280 1457 1300 1477
rect 1320 1457 1340 1477
rect 1360 1457 1380 1477
rect 1400 1457 1420 1477
rect 1440 1457 1460 1477
rect 10 1415 30 1435
rect 50 1415 70 1435
rect 90 1415 110 1435
rect 130 1415 150 1435
rect 1760 1375 1780 1395
rect 1800 1375 1820 1395
rect 1840 1375 1860 1395
rect 1880 1375 1900 1395
rect 1920 1375 1940 1395
rect 1960 1375 1980 1395
rect 2000 1375 2020 1395
rect 2040 1375 2060 1395
rect 2080 1375 2100 1395
rect 2120 1375 2140 1395
rect 2160 1375 2180 1395
rect 2200 1375 2220 1395
rect 2240 1375 2260 1395
rect 2280 1375 2300 1395
rect 2320 1375 2340 1395
rect 2360 1375 2380 1395
rect 2400 1375 2420 1395
rect 2440 1375 2460 1395
rect 2480 1375 2500 1395
rect 2520 1375 2540 1395
rect 10 1335 30 1355
rect 50 1335 70 1355
rect 90 1335 110 1355
rect 130 1335 150 1355
rect 680 1293 700 1313
rect 720 1293 740 1313
rect 760 1293 780 1313
rect 800 1293 820 1313
rect 840 1293 860 1313
rect 880 1293 900 1313
rect 920 1293 940 1313
rect 960 1293 980 1313
rect 1000 1293 1020 1313
rect 1040 1293 1060 1313
rect 1080 1293 1100 1313
rect 1120 1293 1140 1313
rect 1160 1293 1180 1313
rect 1200 1293 1220 1313
rect 1240 1293 1260 1313
rect 1280 1293 1300 1313
rect 1320 1293 1340 1313
rect 1360 1293 1380 1313
rect 1400 1293 1420 1313
rect 1440 1293 1460 1313
rect 10 1250 30 1270
rect 50 1250 70 1270
rect 90 1250 110 1270
rect 130 1250 150 1270
rect 1760 1211 1780 1231
rect 1800 1211 1820 1231
rect 1840 1211 1860 1231
rect 1880 1211 1900 1231
rect 1920 1211 1940 1231
rect 1960 1211 1980 1231
rect 2000 1211 2020 1231
rect 2040 1211 2060 1231
rect 2080 1211 2100 1231
rect 2120 1211 2140 1231
rect 2160 1211 2180 1231
rect 2200 1211 2220 1231
rect 2240 1211 2260 1231
rect 2280 1211 2300 1231
rect 2320 1211 2340 1231
rect 2360 1211 2380 1231
rect 2400 1211 2420 1231
rect 2440 1211 2460 1231
rect 2480 1211 2500 1231
rect 2520 1211 2540 1231
rect 10 1170 30 1190
rect 50 1170 70 1190
rect 90 1170 110 1190
rect 130 1170 150 1190
rect 680 1129 700 1149
rect 720 1129 740 1149
rect 760 1129 780 1149
rect 800 1129 820 1149
rect 840 1129 860 1149
rect 880 1129 900 1149
rect 920 1129 940 1149
rect 960 1129 980 1149
rect 1000 1129 1020 1149
rect 1040 1129 1060 1149
rect 1080 1129 1100 1149
rect 1120 1129 1140 1149
rect 1160 1129 1180 1149
rect 1200 1129 1220 1149
rect 1240 1129 1260 1149
rect 1280 1129 1300 1149
rect 1320 1129 1340 1149
rect 1360 1129 1380 1149
rect 1400 1129 1420 1149
rect 1440 1129 1460 1149
rect 10 1090 30 1110
rect 50 1090 70 1110
rect 90 1090 110 1110
rect 130 1090 150 1110
rect 1760 1047 1780 1067
rect 1800 1047 1820 1067
rect 1840 1047 1860 1067
rect 1880 1047 1900 1067
rect 1920 1047 1940 1067
rect 1960 1047 1980 1067
rect 2000 1047 2020 1067
rect 2040 1047 2060 1067
rect 2080 1047 2100 1067
rect 2120 1047 2140 1067
rect 2160 1047 2180 1067
rect 2200 1047 2220 1067
rect 2240 1047 2260 1067
rect 2280 1047 2300 1067
rect 2320 1047 2340 1067
rect 2360 1047 2380 1067
rect 2400 1047 2420 1067
rect 2440 1047 2460 1067
rect 2480 1047 2500 1067
rect 2520 1047 2540 1067
rect 10 1005 30 1025
rect 50 1005 70 1025
rect 90 1005 110 1025
rect 130 1005 150 1025
rect 680 965 700 985
rect 720 965 740 985
rect 760 965 780 985
rect 800 965 820 985
rect 840 965 860 985
rect 880 965 900 985
rect 920 965 940 985
rect 960 965 980 985
rect 1000 965 1020 985
rect 1040 965 1060 985
rect 1080 965 1100 985
rect 1120 965 1140 985
rect 1160 965 1180 985
rect 1200 965 1220 985
rect 1240 965 1260 985
rect 1280 965 1300 985
rect 1320 965 1340 985
rect 1360 965 1380 985
rect 1400 965 1420 985
rect 1440 965 1460 985
rect 10 925 30 945
rect 50 925 70 945
rect 90 925 110 945
rect 130 925 150 945
rect 1760 883 1780 903
rect 1800 883 1820 903
rect 1840 883 1860 903
rect 1880 883 1900 903
rect 1920 883 1940 903
rect 1960 883 1980 903
rect 2000 883 2020 903
rect 2040 883 2060 903
rect 2080 883 2100 903
rect 2120 883 2140 903
rect 2160 883 2180 903
rect 2200 883 2220 903
rect 2240 883 2260 903
rect 2280 883 2300 903
rect 2320 883 2340 903
rect 2360 883 2380 903
rect 2400 883 2420 903
rect 2440 883 2460 903
rect 2480 883 2500 903
rect 2520 883 2540 903
rect 10 840 30 860
rect 50 840 70 860
rect 90 840 110 860
rect 130 840 150 860
rect 680 801 700 821
rect 720 801 740 821
rect 760 801 780 821
rect 800 801 820 821
rect 840 801 860 821
rect 880 801 900 821
rect 920 801 940 821
rect 960 801 980 821
rect 1000 801 1020 821
rect 1040 801 1060 821
rect 1080 801 1100 821
rect 1120 801 1140 821
rect 1160 801 1180 821
rect 1200 801 1220 821
rect 1240 801 1260 821
rect 1280 801 1300 821
rect 1320 801 1340 821
rect 1360 801 1380 821
rect 1400 801 1420 821
rect 1440 801 1460 821
rect 10 760 30 780
rect 50 760 70 780
rect 90 760 110 780
rect 130 760 150 780
rect 1760 719 1780 739
rect 1800 719 1820 739
rect 1840 719 1860 739
rect 1880 719 1900 739
rect 1920 719 1940 739
rect 1960 719 1980 739
rect 2000 719 2020 739
rect 2040 719 2060 739
rect 2080 719 2100 739
rect 2120 719 2140 739
rect 2160 719 2180 739
rect 2200 719 2220 739
rect 2240 719 2260 739
rect 2280 719 2300 739
rect 2320 719 2340 739
rect 2360 719 2380 739
rect 2400 719 2420 739
rect 2440 719 2460 739
rect 2480 719 2500 739
rect 2520 719 2540 739
rect 10 680 30 700
rect 50 680 70 700
rect 90 680 110 700
rect 130 680 150 700
rect 680 637 700 657
rect 720 637 740 657
rect 760 637 780 657
rect 800 637 820 657
rect 840 637 860 657
rect 880 637 900 657
rect 920 637 940 657
rect 960 637 980 657
rect 1000 637 1020 657
rect 1040 637 1060 657
rect 1080 637 1100 657
rect 1120 637 1140 657
rect 1160 637 1180 657
rect 1200 637 1220 657
rect 1240 637 1260 657
rect 1280 637 1300 657
rect 1320 637 1340 657
rect 1360 637 1380 657
rect 1400 637 1420 657
rect 1440 637 1460 657
rect 10 595 30 615
rect 50 595 70 615
rect 90 595 110 615
rect 130 595 150 615
rect 1760 555 1780 575
rect 1800 555 1820 575
rect 1840 555 1860 575
rect 1880 555 1900 575
rect 1920 555 1940 575
rect 1960 555 1980 575
rect 2000 555 2020 575
rect 2040 555 2060 575
rect 2080 555 2100 575
rect 2120 555 2140 575
rect 2160 555 2180 575
rect 2200 555 2220 575
rect 2240 555 2260 575
rect 2280 555 2300 575
rect 2320 555 2340 575
rect 2360 555 2380 575
rect 2400 555 2420 575
rect 2440 555 2460 575
rect 2480 555 2500 575
rect 2520 555 2540 575
rect 10 515 30 535
rect 50 515 70 535
rect 90 515 110 535
rect 130 515 150 535
rect 680 473 700 493
rect 720 473 740 493
rect 760 473 780 493
rect 800 473 820 493
rect 840 473 860 493
rect 880 473 900 493
rect 920 473 940 493
rect 960 473 980 493
rect 1000 473 1020 493
rect 1040 473 1060 493
rect 1080 473 1100 493
rect 1120 473 1140 493
rect 1160 473 1180 493
rect 1200 473 1220 493
rect 1240 473 1260 493
rect 1280 473 1300 493
rect 1320 473 1340 493
rect 1360 473 1380 493
rect 1400 473 1420 493
rect 1440 473 1460 493
rect 10 435 30 455
rect 50 435 70 455
rect 90 435 110 455
rect 130 435 150 455
rect 1760 391 1780 411
rect 1800 391 1820 411
rect 1840 391 1860 411
rect 1880 391 1900 411
rect 1920 391 1940 411
rect 1960 391 1980 411
rect 2000 391 2020 411
rect 2040 391 2060 411
rect 2080 391 2100 411
rect 2120 391 2140 411
rect 2160 391 2180 411
rect 2200 391 2220 411
rect 2240 391 2260 411
rect 2280 391 2300 411
rect 2320 391 2340 411
rect 2360 391 2380 411
rect 2400 391 2420 411
rect 2440 391 2460 411
rect 2480 391 2500 411
rect 2520 391 2540 411
rect 10 350 30 370
rect 50 350 70 370
rect 90 350 110 370
rect 130 350 150 370
rect 680 309 700 329
rect 720 309 740 329
rect 760 309 780 329
rect 800 309 820 329
rect 840 309 860 329
rect 880 309 900 329
rect 920 309 940 329
rect 960 309 980 329
rect 1000 309 1020 329
rect 1040 309 1060 329
rect 1080 309 1100 329
rect 1120 309 1140 329
rect 1160 309 1180 329
rect 1200 309 1220 329
rect 1240 309 1260 329
rect 1280 309 1300 329
rect 1320 309 1340 329
rect 1360 309 1380 329
rect 1400 309 1420 329
rect 1440 309 1460 329
rect 10 270 30 290
rect 50 270 70 290
rect 90 270 110 290
rect 130 270 150 290
rect 1760 227 1780 247
rect 1800 227 1820 247
rect 1840 227 1860 247
rect 1880 227 1900 247
rect 1920 227 1940 247
rect 1960 227 1980 247
rect 2000 227 2020 247
rect 2040 227 2060 247
rect 2080 227 2100 247
rect 2120 227 2140 247
rect 2160 227 2180 247
rect 2200 227 2220 247
rect 2240 227 2260 247
rect 2280 227 2300 247
rect 2320 227 2340 247
rect 2360 227 2380 247
rect 2400 227 2420 247
rect 2440 227 2460 247
rect 2480 227 2500 247
rect 2520 227 2540 247
rect 10 190 30 210
rect 50 190 70 210
rect 90 190 110 210
rect 130 190 150 210
rect 680 145 700 165
rect 720 145 740 165
rect 760 145 780 165
rect 800 145 820 165
rect 840 145 860 165
rect 880 145 900 165
rect 920 145 940 165
rect 960 145 980 165
rect 1000 145 1020 165
rect 1040 145 1060 165
rect 1080 145 1100 165
rect 1120 145 1140 165
rect 1160 145 1180 165
rect 1200 145 1220 165
rect 1240 145 1260 165
rect 1280 145 1300 165
rect 1320 145 1340 165
rect 1360 145 1380 165
rect 1400 145 1420 165
rect 1440 145 1460 165
rect 320 75 340 95
rect 360 75 380 95
rect 400 75 420 95
rect 1760 75 1780 95
rect 1800 75 1820 95
rect 1840 75 1860 95
rect 1880 75 1900 95
rect 1920 75 1940 95
rect 1960 75 1980 95
rect 2000 75 2020 95
rect 2040 75 2060 95
rect 2080 75 2100 95
rect 2120 75 2140 95
rect 2160 75 2180 95
rect 2200 75 2220 95
rect 2240 75 2260 95
rect 2280 75 2300 95
rect 2320 75 2340 95
rect 2360 75 2380 95
rect 2400 75 2420 95
rect 2440 75 2460 95
rect 2480 75 2500 95
rect 2520 75 2540 95
rect 2560 75 2580 95
rect 2600 75 2620 95
rect 2640 75 2660 95
rect 1760 -30 1780 -10
rect 1800 -30 1820 -10
rect 1840 -30 1860 -10
rect 1880 -30 1900 -10
rect 1920 -30 1940 -10
rect 1960 -30 1980 -10
rect 2000 -30 2020 -10
rect 2040 -30 2060 -10
rect 2080 -30 2100 -10
rect 2120 -30 2140 -10
rect 2160 -30 2180 -10
rect 2200 -30 2220 -10
rect 2240 -30 2260 -10
rect 2280 -30 2300 -10
rect 2320 -30 2340 -10
rect 2360 -30 2380 -10
rect 2400 -30 2420 -10
rect 2440 -30 2460 -10
rect 2480 -30 2500 -10
rect 2520 -30 2540 -10
rect 1760 -70 1780 -50
rect 1800 -70 1820 -50
rect 1840 -70 1860 -50
rect 1880 -70 1900 -50
rect 1920 -70 1940 -50
rect 1960 -70 1980 -50
rect 2000 -70 2020 -50
rect 2040 -70 2060 -50
rect 2080 -70 2100 -50
rect 2120 -70 2140 -50
rect 2160 -70 2180 -50
rect 2200 -70 2220 -50
rect 2240 -70 2260 -50
rect 2280 -70 2300 -50
rect 2320 -70 2340 -50
rect 2360 -70 2380 -50
rect 2400 -70 2420 -50
rect 2440 -70 2460 -50
rect 2480 -70 2500 -50
rect 2520 -70 2540 -50
rect -60 -120 -40 -95
rect -20 -120 0 -95
rect 20 -120 40 -95
rect 60 -120 80 -95
rect 680 -165 700 -145
rect 720 -165 740 -145
rect 760 -165 780 -145
rect 800 -165 820 -145
rect 840 -165 860 -145
rect 880 -165 900 -145
rect 920 -165 940 -145
rect 960 -165 980 -145
rect 1000 -165 1020 -145
rect 1040 -165 1060 -145
rect 1080 -165 1100 -145
rect 1120 -165 1140 -145
rect 1160 -165 1180 -145
rect 1200 -165 1220 -145
rect 1240 -165 1260 -145
rect 1280 -165 1300 -145
rect 1320 -165 1340 -145
rect 1360 -165 1380 -145
rect 1400 -165 1420 -145
rect 1440 -165 1460 -145
rect -60 -215 -40 -190
rect -20 -215 0 -190
rect 20 -215 40 -190
rect 60 -215 80 -190
rect 1760 -260 1780 -240
rect 1800 -260 1820 -240
rect 1840 -260 1860 -240
rect 1880 -260 1900 -240
rect 1920 -260 1940 -240
rect 1960 -260 1980 -240
rect 2000 -260 2020 -240
rect 2040 -260 2060 -240
rect 2080 -260 2100 -240
rect 2120 -260 2140 -240
rect 2160 -260 2180 -240
rect 2200 -260 2220 -240
rect 2240 -260 2260 -240
rect 2280 -260 2300 -240
rect 2320 -260 2340 -240
rect 2360 -260 2380 -240
rect 2400 -260 2420 -240
rect 2440 -260 2460 -240
rect 2480 -260 2500 -240
rect 2520 -260 2540 -240
rect -60 -310 -40 -285
rect -20 -310 0 -285
rect 20 -310 40 -285
rect 60 -310 80 -285
rect 680 -355 700 -335
rect 720 -355 740 -335
rect 760 -355 780 -335
rect 800 -355 820 -335
rect 840 -355 860 -335
rect 880 -355 900 -335
rect 920 -355 940 -335
rect 960 -355 980 -335
rect 1000 -355 1020 -335
rect 1040 -355 1060 -335
rect 1080 -355 1100 -335
rect 1120 -355 1140 -335
rect 1160 -355 1180 -335
rect 1200 -355 1220 -335
rect 1240 -355 1260 -335
rect 1280 -355 1300 -335
rect 1320 -355 1340 -335
rect 1360 -355 1380 -335
rect 1400 -355 1420 -335
rect 1440 -355 1460 -335
rect -60 -405 -40 -380
rect -20 -405 0 -380
rect 20 -405 40 -380
rect 60 -405 80 -380
rect 1760 -450 1780 -430
rect 1800 -450 1820 -430
rect 1840 -450 1860 -430
rect 1880 -450 1900 -430
rect 1920 -450 1940 -430
rect 1960 -450 1980 -430
rect 2000 -450 2020 -430
rect 2040 -450 2060 -430
rect 2080 -450 2100 -430
rect 2120 -450 2140 -430
rect 2160 -450 2180 -430
rect 2200 -450 2220 -430
rect 2240 -450 2260 -430
rect 2280 -450 2300 -430
rect 2320 -450 2340 -430
rect 2360 -450 2380 -430
rect 2400 -450 2420 -430
rect 2440 -450 2460 -430
rect 2480 -450 2500 -430
rect 2520 -450 2540 -430
rect -60 -500 -40 -475
rect -20 -500 0 -475
rect 20 -500 40 -475
rect 60 -500 80 -475
rect 680 -545 700 -525
rect 720 -545 740 -525
rect 760 -545 780 -525
rect 800 -545 820 -525
rect 840 -545 860 -525
rect 880 -545 900 -525
rect 920 -545 940 -525
rect 960 -545 980 -525
rect 1000 -545 1020 -525
rect 1040 -545 1060 -525
rect 1080 -545 1100 -525
rect 1120 -545 1140 -525
rect 1160 -545 1180 -525
rect 1200 -545 1220 -525
rect 1240 -545 1260 -525
rect 1280 -545 1300 -525
rect 1320 -545 1340 -525
rect 1360 -545 1380 -525
rect 1400 -545 1420 -525
rect 1440 -545 1460 -525
rect -60 -595 -40 -570
rect -20 -595 0 -570
rect 20 -595 40 -570
rect 60 -595 80 -570
rect 1760 -640 1780 -620
rect 1800 -640 1820 -620
rect 1840 -640 1860 -620
rect 1880 -640 1900 -620
rect 1920 -640 1940 -620
rect 1960 -640 1980 -620
rect 2000 -640 2020 -620
rect 2040 -640 2060 -620
rect 2080 -640 2100 -620
rect 2120 -640 2140 -620
rect 2160 -640 2180 -620
rect 2200 -640 2220 -620
rect 2240 -640 2260 -620
rect 2280 -640 2300 -620
rect 2320 -640 2340 -620
rect 2360 -640 2380 -620
rect 2400 -640 2420 -620
rect 2440 -640 2460 -620
rect 2480 -640 2500 -620
rect 2520 -640 2540 -620
rect -60 -690 -40 -665
rect -20 -690 0 -665
rect 20 -690 40 -665
rect 60 -690 80 -665
rect 680 -735 700 -715
rect 720 -735 740 -715
rect 760 -735 780 -715
rect 800 -735 820 -715
rect 840 -735 860 -715
rect 880 -735 900 -715
rect 920 -735 940 -715
rect 960 -735 980 -715
rect 1000 -735 1020 -715
rect 1040 -735 1060 -715
rect 1080 -735 1100 -715
rect 1120 -735 1140 -715
rect 1160 -735 1180 -715
rect 1200 -735 1220 -715
rect 1240 -735 1260 -715
rect 1280 -735 1300 -715
rect 1320 -735 1340 -715
rect 1360 -735 1380 -715
rect 1400 -735 1420 -715
rect 1440 -735 1460 -715
rect -60 -785 -40 -760
rect -20 -785 0 -760
rect 20 -785 40 -760
rect 60 -785 80 -760
rect 1760 -830 1780 -810
rect 1800 -830 1820 -810
rect 1840 -830 1860 -810
rect 1880 -830 1900 -810
rect 1920 -830 1940 -810
rect 1960 -830 1980 -810
rect 2000 -830 2020 -810
rect 2040 -830 2060 -810
rect 2080 -830 2100 -810
rect 2120 -830 2140 -810
rect 2160 -830 2180 -810
rect 2200 -830 2220 -810
rect 2240 -830 2260 -810
rect 2280 -830 2300 -810
rect 2320 -830 2340 -810
rect 2360 -830 2380 -810
rect 2400 -830 2420 -810
rect 2440 -830 2460 -810
rect 2480 -830 2500 -810
rect 2520 -830 2540 -810
rect -60 -880 -40 -855
rect -20 -880 0 -855
rect 20 -880 40 -855
rect 60 -880 80 -855
rect 680 -925 700 -905
rect 720 -925 740 -905
rect 760 -925 780 -905
rect 800 -925 820 -905
rect 840 -925 860 -905
rect 880 -925 900 -905
rect 920 -925 940 -905
rect 960 -925 980 -905
rect 1000 -925 1020 -905
rect 1040 -925 1060 -905
rect 1080 -925 1100 -905
rect 1120 -925 1140 -905
rect 1160 -925 1180 -905
rect 1200 -925 1220 -905
rect 1240 -925 1260 -905
rect 1280 -925 1300 -905
rect 1320 -925 1340 -905
rect 1360 -925 1380 -905
rect 1400 -925 1420 -905
rect 1440 -925 1460 -905
rect -60 -975 -40 -950
rect -20 -975 0 -950
rect 20 -975 40 -950
rect 60 -975 80 -950
rect 1760 -1020 1780 -1000
rect 1800 -1020 1820 -1000
rect 1840 -1020 1860 -1000
rect 1880 -1020 1900 -1000
rect 1920 -1020 1940 -1000
rect 1960 -1020 1980 -1000
rect 2000 -1020 2020 -1000
rect 2040 -1020 2060 -1000
rect 2080 -1020 2100 -1000
rect 2120 -1020 2140 -1000
rect 2160 -1020 2180 -1000
rect 2200 -1020 2220 -1000
rect 2240 -1020 2260 -1000
rect 2280 -1020 2300 -1000
rect 2320 -1020 2340 -1000
rect 2360 -1020 2380 -1000
rect 2400 -1020 2420 -1000
rect 2440 -1020 2460 -1000
rect 2480 -1020 2500 -1000
rect 2520 -1020 2540 -1000
rect -60 -1070 -40 -1045
rect -20 -1070 0 -1045
rect 20 -1070 40 -1045
rect 60 -1070 80 -1045
rect 680 -1115 700 -1095
rect 720 -1115 740 -1095
rect 760 -1115 780 -1095
rect 800 -1115 820 -1095
rect 840 -1115 860 -1095
rect 880 -1115 900 -1095
rect 920 -1115 940 -1095
rect 960 -1115 980 -1095
rect 1000 -1115 1020 -1095
rect 1040 -1115 1060 -1095
rect 1080 -1115 1100 -1095
rect 1120 -1115 1140 -1095
rect 1160 -1115 1180 -1095
rect 1200 -1115 1220 -1095
rect 1240 -1115 1260 -1095
rect 1280 -1115 1300 -1095
rect 1320 -1115 1340 -1095
rect 1360 -1115 1380 -1095
rect 1400 -1115 1420 -1095
rect 1440 -1115 1460 -1095
rect -60 -1165 -40 -1140
rect -20 -1165 0 -1140
rect 20 -1165 40 -1140
rect 60 -1165 80 -1140
rect 1760 -1210 1780 -1190
rect 1800 -1210 1820 -1190
rect 1840 -1210 1860 -1190
rect 1880 -1210 1900 -1190
rect 1920 -1210 1940 -1190
rect 1960 -1210 1980 -1190
rect 2000 -1210 2020 -1190
rect 2040 -1210 2060 -1190
rect 2080 -1210 2100 -1190
rect 2120 -1210 2140 -1190
rect 2160 -1210 2180 -1190
rect 2200 -1210 2220 -1190
rect 2240 -1210 2260 -1190
rect 2280 -1210 2300 -1190
rect 2320 -1210 2340 -1190
rect 2360 -1210 2380 -1190
rect 2400 -1210 2420 -1190
rect 2440 -1210 2460 -1190
rect 2480 -1210 2500 -1190
rect 2520 -1210 2540 -1190
rect -60 -1260 -40 -1235
rect -20 -1260 0 -1235
rect 20 -1260 40 -1235
rect 60 -1260 80 -1235
rect 680 -1305 700 -1285
rect 720 -1305 740 -1285
rect 760 -1305 780 -1285
rect 800 -1305 820 -1285
rect 840 -1305 860 -1285
rect 880 -1305 900 -1285
rect 920 -1305 940 -1285
rect 960 -1305 980 -1285
rect 1000 -1305 1020 -1285
rect 1040 -1305 1060 -1285
rect 1080 -1305 1100 -1285
rect 1120 -1305 1140 -1285
rect 1160 -1305 1180 -1285
rect 1200 -1305 1220 -1285
rect 1240 -1305 1260 -1285
rect 1280 -1305 1300 -1285
rect 1320 -1305 1340 -1285
rect 1360 -1305 1380 -1285
rect 1400 -1305 1420 -1285
rect 1440 -1305 1460 -1285
rect -60 -1355 -40 -1330
rect -20 -1355 0 -1330
rect 20 -1355 40 -1330
rect 60 -1355 80 -1330
rect 1760 -1400 1780 -1380
rect 1800 -1400 1820 -1380
rect 1840 -1400 1860 -1380
rect 1880 -1400 1900 -1380
rect 1920 -1400 1940 -1380
rect 1960 -1400 1980 -1380
rect 2000 -1400 2020 -1380
rect 2040 -1400 2060 -1380
rect 2080 -1400 2100 -1380
rect 2120 -1400 2140 -1380
rect 2160 -1400 2180 -1380
rect 2200 -1400 2220 -1380
rect 2240 -1400 2260 -1380
rect 2280 -1400 2300 -1380
rect 2320 -1400 2340 -1380
rect 2360 -1400 2380 -1380
rect 2400 -1400 2420 -1380
rect 2440 -1400 2460 -1380
rect 2480 -1400 2500 -1380
rect 2520 -1400 2540 -1380
rect -60 -1450 -40 -1425
rect -20 -1450 0 -1425
rect 20 -1450 40 -1425
rect 60 -1450 80 -1425
rect 680 -1495 700 -1475
rect 720 -1495 740 -1475
rect 760 -1495 780 -1475
rect 800 -1495 820 -1475
rect 840 -1495 860 -1475
rect 880 -1495 900 -1475
rect 920 -1495 940 -1475
rect 960 -1495 980 -1475
rect 1000 -1495 1020 -1475
rect 1040 -1495 1060 -1475
rect 1080 -1495 1100 -1475
rect 1120 -1495 1140 -1475
rect 1160 -1495 1180 -1475
rect 1200 -1495 1220 -1475
rect 1240 -1495 1260 -1475
rect 1280 -1495 1300 -1475
rect 1320 -1495 1340 -1475
rect 1360 -1495 1380 -1475
rect 1400 -1495 1420 -1475
rect 1440 -1495 1460 -1475
rect -60 -1545 -40 -1520
rect -20 -1545 0 -1520
rect 20 -1545 40 -1520
rect 60 -1545 80 -1520
rect 1760 -1590 1780 -1570
rect 1800 -1590 1820 -1570
rect 1840 -1590 1860 -1570
rect 1880 -1590 1900 -1570
rect 1920 -1590 1940 -1570
rect 1960 -1590 1980 -1570
rect 2000 -1590 2020 -1570
rect 2040 -1590 2060 -1570
rect 2080 -1590 2100 -1570
rect 2120 -1590 2140 -1570
rect 2160 -1590 2180 -1570
rect 2200 -1590 2220 -1570
rect 2240 -1590 2260 -1570
rect 2280 -1590 2300 -1570
rect 2320 -1590 2340 -1570
rect 2360 -1590 2380 -1570
rect 2400 -1590 2420 -1570
rect 2440 -1590 2460 -1570
rect 2480 -1590 2500 -1570
rect 2520 -1590 2540 -1570
rect -60 -1640 -40 -1615
rect -20 -1640 0 -1615
rect 20 -1640 40 -1615
rect 60 -1640 80 -1615
rect 680 -1685 700 -1665
rect 720 -1685 740 -1665
rect 760 -1685 780 -1665
rect 800 -1685 820 -1665
rect 840 -1685 860 -1665
rect 880 -1685 900 -1665
rect 920 -1685 940 -1665
rect 960 -1685 980 -1665
rect 1000 -1685 1020 -1665
rect 1040 -1685 1060 -1665
rect 1080 -1685 1100 -1665
rect 1120 -1685 1140 -1665
rect 1160 -1685 1180 -1665
rect 1200 -1685 1220 -1665
rect 1240 -1685 1260 -1665
rect 1280 -1685 1300 -1665
rect 1320 -1685 1340 -1665
rect 1360 -1685 1380 -1665
rect 1400 -1685 1420 -1665
rect 1440 -1685 1460 -1665
rect -60 -1735 -40 -1710
rect -20 -1735 0 -1710
rect 20 -1735 40 -1710
rect 60 -1735 80 -1710
rect 1760 -1780 1780 -1760
rect 1800 -1780 1820 -1760
rect 1840 -1780 1860 -1760
rect 1880 -1780 1900 -1760
rect 1920 -1780 1940 -1760
rect 1960 -1780 1980 -1760
rect 2000 -1780 2020 -1760
rect 2040 -1780 2060 -1760
rect 2080 -1780 2100 -1760
rect 2120 -1780 2140 -1760
rect 2160 -1780 2180 -1760
rect 2200 -1780 2220 -1760
rect 2240 -1780 2260 -1760
rect 2280 -1780 2300 -1760
rect 2320 -1780 2340 -1760
rect 2360 -1780 2380 -1760
rect 2400 -1780 2420 -1760
rect 2440 -1780 2460 -1760
rect 2480 -1780 2500 -1760
rect 2520 -1780 2540 -1760
rect -60 -1830 -40 -1805
rect -20 -1830 0 -1805
rect 20 -1830 40 -1805
rect 60 -1830 80 -1805
rect 680 -1875 700 -1855
rect 720 -1875 740 -1855
rect 760 -1875 780 -1855
rect 800 -1875 820 -1855
rect 840 -1875 860 -1855
rect 880 -1875 900 -1855
rect 920 -1875 940 -1855
rect 960 -1875 980 -1855
rect 1000 -1875 1020 -1855
rect 1040 -1875 1060 -1855
rect 1080 -1875 1100 -1855
rect 1120 -1875 1140 -1855
rect 1160 -1875 1180 -1855
rect 1200 -1875 1220 -1855
rect 1240 -1875 1260 -1855
rect 1280 -1875 1300 -1855
rect 1320 -1875 1340 -1855
rect 1360 -1875 1380 -1855
rect 1400 -1875 1420 -1855
rect 1440 -1875 1460 -1855
rect -60 -1925 -40 -1900
rect -20 -1925 0 -1900
rect 20 -1925 40 -1900
rect 60 -1925 80 -1900
rect 1760 -1970 1780 -1950
rect 1800 -1970 1820 -1950
rect 1840 -1970 1860 -1950
rect 1880 -1970 1900 -1950
rect 1920 -1970 1940 -1950
rect 1960 -1970 1980 -1950
rect 2000 -1970 2020 -1950
rect 2040 -1970 2060 -1950
rect 2080 -1970 2100 -1950
rect 2120 -1970 2140 -1950
rect 2160 -1970 2180 -1950
rect 2200 -1970 2220 -1950
rect 2240 -1970 2260 -1950
rect 2280 -1970 2300 -1950
rect 2320 -1970 2340 -1950
rect 2360 -1970 2380 -1950
rect 2400 -1970 2420 -1950
rect 2440 -1970 2460 -1950
rect 2480 -1970 2500 -1950
rect 2520 -1970 2540 -1950
rect -60 -2020 -40 -1995
rect -20 -2020 0 -1995
rect 20 -2020 40 -1995
rect 60 -2020 80 -1995
rect 680 -2065 700 -2045
rect 720 -2065 740 -2045
rect 760 -2065 780 -2045
rect 800 -2065 820 -2045
rect 840 -2065 860 -2045
rect 880 -2065 900 -2045
rect 920 -2065 940 -2045
rect 960 -2065 980 -2045
rect 1000 -2065 1020 -2045
rect 1040 -2065 1060 -2045
rect 1080 -2065 1100 -2045
rect 1120 -2065 1140 -2045
rect 1160 -2065 1180 -2045
rect 1200 -2065 1220 -2045
rect 1240 -2065 1260 -2045
rect 1280 -2065 1300 -2045
rect 1320 -2065 1340 -2045
rect 1360 -2065 1380 -2045
rect 1400 -2065 1420 -2045
rect 1440 -2065 1460 -2045
rect -60 -2115 -40 -2090
rect -20 -2115 0 -2090
rect 20 -2115 40 -2090
rect 60 -2115 80 -2090
rect 1760 -2160 1780 -2140
rect 1800 -2160 1820 -2140
rect 1840 -2160 1860 -2140
rect 1880 -2160 1900 -2140
rect 1920 -2160 1940 -2140
rect 1960 -2160 1980 -2140
rect 2000 -2160 2020 -2140
rect 2040 -2160 2060 -2140
rect 2080 -2160 2100 -2140
rect 2120 -2160 2140 -2140
rect 2160 -2160 2180 -2140
rect 2200 -2160 2220 -2140
rect 2240 -2160 2260 -2140
rect 2280 -2160 2300 -2140
rect 2320 -2160 2340 -2140
rect 2360 -2160 2380 -2140
rect 2400 -2160 2420 -2140
rect 2440 -2160 2460 -2140
rect 2480 -2160 2500 -2140
rect 2520 -2160 2540 -2140
rect -60 -2210 -40 -2185
rect -20 -2210 0 -2185
rect 20 -2210 40 -2185
rect 60 -2210 80 -2185
rect 680 -2255 700 -2235
rect 720 -2255 740 -2235
rect 760 -2255 780 -2235
rect 800 -2255 820 -2235
rect 840 -2255 860 -2235
rect 880 -2255 900 -2235
rect 920 -2255 940 -2235
rect 960 -2255 980 -2235
rect 1000 -2255 1020 -2235
rect 1040 -2255 1060 -2235
rect 1080 -2255 1100 -2235
rect 1120 -2255 1140 -2235
rect 1160 -2255 1180 -2235
rect 1200 -2255 1220 -2235
rect 1240 -2255 1260 -2235
rect 1280 -2255 1300 -2235
rect 1320 -2255 1340 -2235
rect 1360 -2255 1380 -2235
rect 1400 -2255 1420 -2235
rect 1440 -2255 1460 -2235
rect -60 -2305 -40 -2280
rect -20 -2305 0 -2280
rect 20 -2305 40 -2280
rect 60 -2305 80 -2280
rect 1760 -2350 1780 -2330
rect 1800 -2350 1820 -2330
rect 1840 -2350 1860 -2330
rect 1880 -2350 1900 -2330
rect 1920 -2350 1940 -2330
rect 1960 -2350 1980 -2330
rect 2000 -2350 2020 -2330
rect 2040 -2350 2060 -2330
rect 2080 -2350 2100 -2330
rect 2120 -2350 2140 -2330
rect 2160 -2350 2180 -2330
rect 2200 -2350 2220 -2330
rect 2240 -2350 2260 -2330
rect 2280 -2350 2300 -2330
rect 2320 -2350 2340 -2330
rect 2360 -2350 2380 -2330
rect 2400 -2350 2420 -2330
rect 2440 -2350 2460 -2330
rect 2480 -2350 2500 -2330
rect 2520 -2350 2540 -2330
rect -60 -2400 -40 -2375
rect -20 -2400 0 -2375
rect 20 -2400 40 -2375
rect 60 -2400 80 -2375
rect 680 -2445 700 -2425
rect 720 -2445 740 -2425
rect 760 -2445 780 -2425
rect 800 -2445 820 -2425
rect 840 -2445 860 -2425
rect 880 -2445 900 -2425
rect 920 -2445 940 -2425
rect 960 -2445 980 -2425
rect 1000 -2445 1020 -2425
rect 1040 -2445 1060 -2425
rect 1080 -2445 1100 -2425
rect 1120 -2445 1140 -2425
rect 1160 -2445 1180 -2425
rect 1200 -2445 1220 -2425
rect 1240 -2445 1260 -2425
rect 1280 -2445 1300 -2425
rect 1320 -2445 1340 -2425
rect 1360 -2445 1380 -2425
rect 1400 -2445 1420 -2425
rect 1440 -2445 1460 -2425
rect -60 -2495 -40 -2470
rect -20 -2495 0 -2470
rect 20 -2495 40 -2470
rect 60 -2495 80 -2470
rect 1760 -2540 1780 -2520
rect 1800 -2540 1820 -2520
rect 1840 -2540 1860 -2520
rect 1880 -2540 1900 -2520
rect 1920 -2540 1940 -2520
rect 1960 -2540 1980 -2520
rect 2000 -2540 2020 -2520
rect 2040 -2540 2060 -2520
rect 2080 -2540 2100 -2520
rect 2120 -2540 2140 -2520
rect 2160 -2540 2180 -2520
rect 2200 -2540 2220 -2520
rect 2240 -2540 2260 -2520
rect 2280 -2540 2300 -2520
rect 2320 -2540 2340 -2520
rect 2360 -2540 2380 -2520
rect 2400 -2540 2420 -2520
rect 2440 -2540 2460 -2520
rect 2480 -2540 2500 -2520
rect 2520 -2540 2540 -2520
rect 1760 -2580 1780 -2560
rect 1800 -2580 1820 -2560
rect 1840 -2580 1860 -2560
rect 1880 -2580 1900 -2560
rect 1920 -2580 1940 -2560
rect 1960 -2580 1980 -2560
rect 2000 -2580 2020 -2560
rect 2040 -2580 2060 -2560
rect 2080 -2580 2100 -2560
rect 2120 -2580 2140 -2560
rect 2160 -2580 2180 -2560
rect 2200 -2580 2220 -2560
rect 2240 -2580 2260 -2560
rect 2280 -2580 2300 -2560
rect 2320 -2580 2340 -2560
rect 2360 -2580 2380 -2560
rect 2400 -2580 2420 -2560
rect 2440 -2580 2460 -2560
rect 2480 -2580 2500 -2560
rect 2520 -2580 2540 -2560
<< metal1 >>
rect 175 2365 1070 2375
rect 175 2345 200 2365
rect 220 2345 240 2365
rect 260 2345 280 2365
rect 300 2345 320 2365
rect 340 2345 360 2365
rect 380 2345 400 2365
rect 420 2345 440 2365
rect 460 2345 480 2365
rect 500 2345 520 2365
rect 540 2345 560 2365
rect 580 2345 600 2365
rect 620 2345 640 2365
rect 660 2345 680 2365
rect 700 2345 720 2365
rect 740 2345 760 2365
rect 780 2345 800 2365
rect 820 2345 840 2365
rect 860 2345 880 2365
rect 900 2345 920 2365
rect 940 2345 960 2365
rect 980 2345 1000 2365
rect 1020 2345 1040 2365
rect 1060 2345 1070 2365
rect 175 2335 1070 2345
rect 0 2255 165 2265
rect 0 2235 10 2255
rect 30 2235 50 2255
rect 70 2235 90 2255
rect 110 2235 130 2255
rect 150 2235 165 2255
rect 0 2175 165 2235
rect 0 2155 10 2175
rect 30 2155 50 2175
rect 70 2155 90 2175
rect 110 2155 130 2175
rect 150 2155 165 2175
rect 0 2090 165 2155
rect 0 2070 10 2090
rect 30 2070 50 2090
rect 70 2070 90 2090
rect 110 2070 130 2090
rect 150 2070 165 2090
rect 0 2010 165 2070
rect 0 1990 10 2010
rect 30 1990 50 2010
rect 70 1990 90 2010
rect 110 1990 130 2010
rect 150 1990 165 2010
rect 0 1930 165 1990
rect 0 1910 10 1930
rect 30 1910 50 1930
rect 70 1910 90 1930
rect 110 1910 130 1930
rect 150 1910 165 1930
rect 0 1845 165 1910
rect 0 1825 10 1845
rect 30 1825 50 1845
rect 70 1825 90 1845
rect 110 1825 130 1845
rect 150 1825 165 1845
rect 0 1765 165 1825
rect 0 1745 10 1765
rect 30 1745 50 1765
rect 70 1745 90 1765
rect 110 1745 130 1765
rect 150 1745 165 1765
rect 0 1680 165 1745
rect 0 1660 10 1680
rect 30 1660 50 1680
rect 70 1660 90 1680
rect 110 1660 130 1680
rect 150 1660 165 1680
rect 0 1600 165 1660
rect 0 1580 10 1600
rect 30 1580 50 1600
rect 70 1580 90 1600
rect 110 1580 130 1600
rect 150 1580 165 1600
rect 0 1520 165 1580
rect 0 1500 10 1520
rect 30 1500 50 1520
rect 70 1500 90 1520
rect 110 1500 130 1520
rect 150 1500 165 1520
rect 0 1435 165 1500
rect 0 1415 10 1435
rect 30 1415 50 1435
rect 70 1415 90 1435
rect 110 1415 130 1435
rect 150 1415 165 1435
rect 0 1355 165 1415
rect 0 1335 10 1355
rect 30 1335 50 1355
rect 70 1335 90 1355
rect 110 1335 130 1355
rect 150 1335 165 1355
rect 0 1270 165 1335
rect 0 1250 10 1270
rect 30 1250 50 1270
rect 70 1250 90 1270
rect 110 1250 130 1270
rect 150 1250 165 1270
rect 0 1190 165 1250
rect 0 1170 10 1190
rect 30 1170 50 1190
rect 70 1170 90 1190
rect 110 1170 130 1190
rect 150 1170 165 1190
rect 0 1110 165 1170
rect 0 1090 10 1110
rect 30 1090 50 1110
rect 70 1090 90 1110
rect 110 1090 130 1110
rect 150 1090 165 1110
rect 0 1025 165 1090
rect 0 1005 10 1025
rect 30 1005 50 1025
rect 70 1005 90 1025
rect 110 1005 130 1025
rect 150 1005 165 1025
rect 0 945 165 1005
rect 0 925 10 945
rect 30 925 50 945
rect 70 925 90 945
rect 110 925 130 945
rect 150 925 165 945
rect 0 860 165 925
rect 0 840 10 860
rect 30 840 50 860
rect 70 840 90 860
rect 110 840 130 860
rect 150 840 165 860
rect 0 780 165 840
rect 0 760 10 780
rect 30 760 50 780
rect 70 760 90 780
rect 110 760 130 780
rect 150 760 165 780
rect 0 700 165 760
rect 0 680 10 700
rect 30 680 50 700
rect 70 680 90 700
rect 110 680 130 700
rect 150 680 165 700
rect 0 615 165 680
rect 0 595 10 615
rect 30 595 50 615
rect 70 595 90 615
rect 110 595 130 615
rect 150 595 165 615
rect 0 535 165 595
rect 0 515 10 535
rect 30 515 50 535
rect 70 515 90 535
rect 110 515 130 535
rect 150 515 165 535
rect 0 455 165 515
rect 0 435 10 455
rect 30 435 50 455
rect 70 435 90 455
rect 110 435 130 455
rect 150 435 165 455
rect 0 370 165 435
rect 0 350 10 370
rect 30 350 50 370
rect 70 350 90 370
rect 110 350 130 370
rect 150 350 165 370
rect 0 290 165 350
rect 0 270 10 290
rect 30 270 50 290
rect 70 270 90 290
rect 110 270 130 290
rect 150 270 165 290
rect 0 210 165 270
rect 0 190 10 210
rect 30 190 50 210
rect 70 190 90 210
rect 110 190 130 210
rect 150 190 165 210
rect 0 180 165 190
rect 310 95 430 2335
rect 310 75 320 95
rect 340 75 360 95
rect 380 75 400 95
rect 420 75 430 95
rect 310 65 430 75
rect 670 2297 1470 2307
rect 670 2277 680 2297
rect 700 2277 720 2297
rect 740 2277 760 2297
rect 780 2277 800 2297
rect 820 2277 840 2297
rect 860 2277 880 2297
rect 900 2277 920 2297
rect 940 2277 960 2297
rect 980 2277 1000 2297
rect 1020 2277 1040 2297
rect 1060 2277 1080 2297
rect 1100 2277 1120 2297
rect 1140 2277 1160 2297
rect 1180 2277 1200 2297
rect 1220 2277 1240 2297
rect 1260 2277 1280 2297
rect 1300 2277 1320 2297
rect 1340 2277 1360 2297
rect 1380 2277 1400 2297
rect 1420 2277 1440 2297
rect 1460 2277 1470 2297
rect 670 2133 1470 2277
rect 670 2113 680 2133
rect 700 2113 720 2133
rect 740 2113 760 2133
rect 780 2113 800 2133
rect 820 2113 840 2133
rect 860 2113 880 2133
rect 900 2113 920 2133
rect 940 2113 960 2133
rect 980 2113 1000 2133
rect 1020 2113 1040 2133
rect 1060 2113 1080 2133
rect 1100 2113 1120 2133
rect 1140 2113 1160 2133
rect 1180 2113 1200 2133
rect 1220 2113 1240 2133
rect 1260 2113 1280 2133
rect 1300 2113 1320 2133
rect 1340 2113 1360 2133
rect 1380 2113 1400 2133
rect 1420 2113 1440 2133
rect 1460 2113 1470 2133
rect 670 1969 1470 2113
rect 670 1949 680 1969
rect 700 1949 720 1969
rect 740 1949 760 1969
rect 780 1949 800 1969
rect 820 1949 840 1969
rect 860 1949 880 1969
rect 900 1949 920 1969
rect 940 1949 960 1969
rect 980 1949 1000 1969
rect 1020 1949 1040 1969
rect 1060 1949 1080 1969
rect 1100 1949 1120 1969
rect 1140 1949 1160 1969
rect 1180 1949 1200 1969
rect 1220 1949 1240 1969
rect 1260 1949 1280 1969
rect 1300 1949 1320 1969
rect 1340 1949 1360 1969
rect 1380 1949 1400 1969
rect 1420 1949 1440 1969
rect 1460 1949 1470 1969
rect 670 1805 1470 1949
rect 670 1785 680 1805
rect 700 1785 720 1805
rect 740 1785 760 1805
rect 780 1785 800 1805
rect 820 1785 840 1805
rect 860 1785 880 1805
rect 900 1785 920 1805
rect 940 1785 960 1805
rect 980 1785 1000 1805
rect 1020 1785 1040 1805
rect 1060 1785 1080 1805
rect 1100 1785 1120 1805
rect 1140 1785 1160 1805
rect 1180 1785 1200 1805
rect 1220 1785 1240 1805
rect 1260 1785 1280 1805
rect 1300 1785 1320 1805
rect 1340 1785 1360 1805
rect 1380 1785 1400 1805
rect 1420 1785 1440 1805
rect 1460 1785 1470 1805
rect 670 1641 1470 1785
rect 670 1621 680 1641
rect 700 1621 720 1641
rect 740 1621 760 1641
rect 780 1621 800 1641
rect 820 1621 840 1641
rect 860 1621 880 1641
rect 900 1621 920 1641
rect 940 1621 960 1641
rect 980 1621 1000 1641
rect 1020 1621 1040 1641
rect 1060 1621 1080 1641
rect 1100 1621 1120 1641
rect 1140 1621 1160 1641
rect 1180 1621 1200 1641
rect 1220 1621 1240 1641
rect 1260 1621 1280 1641
rect 1300 1621 1320 1641
rect 1340 1621 1360 1641
rect 1380 1621 1400 1641
rect 1420 1621 1440 1641
rect 1460 1621 1470 1641
rect 670 1477 1470 1621
rect 670 1457 680 1477
rect 700 1457 720 1477
rect 740 1457 760 1477
rect 780 1457 800 1477
rect 820 1457 840 1477
rect 860 1457 880 1477
rect 900 1457 920 1477
rect 940 1457 960 1477
rect 980 1457 1000 1477
rect 1020 1457 1040 1477
rect 1060 1457 1080 1477
rect 1100 1457 1120 1477
rect 1140 1457 1160 1477
rect 1180 1457 1200 1477
rect 1220 1457 1240 1477
rect 1260 1457 1280 1477
rect 1300 1457 1320 1477
rect 1340 1457 1360 1477
rect 1380 1457 1400 1477
rect 1420 1457 1440 1477
rect 1460 1457 1470 1477
rect 670 1313 1470 1457
rect 670 1293 680 1313
rect 700 1293 720 1313
rect 740 1293 760 1313
rect 780 1293 800 1313
rect 820 1293 840 1313
rect 860 1293 880 1313
rect 900 1293 920 1313
rect 940 1293 960 1313
rect 980 1293 1000 1313
rect 1020 1293 1040 1313
rect 1060 1293 1080 1313
rect 1100 1293 1120 1313
rect 1140 1293 1160 1313
rect 1180 1293 1200 1313
rect 1220 1293 1240 1313
rect 1260 1293 1280 1313
rect 1300 1293 1320 1313
rect 1340 1293 1360 1313
rect 1380 1293 1400 1313
rect 1420 1293 1440 1313
rect 1460 1293 1470 1313
rect 670 1149 1470 1293
rect 670 1129 680 1149
rect 700 1129 720 1149
rect 740 1129 760 1149
rect 780 1129 800 1149
rect 820 1129 840 1149
rect 860 1129 880 1149
rect 900 1129 920 1149
rect 940 1129 960 1149
rect 980 1129 1000 1149
rect 1020 1129 1040 1149
rect 1060 1129 1080 1149
rect 1100 1129 1120 1149
rect 1140 1129 1160 1149
rect 1180 1129 1200 1149
rect 1220 1129 1240 1149
rect 1260 1129 1280 1149
rect 1300 1129 1320 1149
rect 1340 1129 1360 1149
rect 1380 1129 1400 1149
rect 1420 1129 1440 1149
rect 1460 1129 1470 1149
rect 670 985 1470 1129
rect 670 965 680 985
rect 700 965 720 985
rect 740 965 760 985
rect 780 965 800 985
rect 820 965 840 985
rect 860 965 880 985
rect 900 965 920 985
rect 940 965 960 985
rect 980 965 1000 985
rect 1020 965 1040 985
rect 1060 965 1080 985
rect 1100 965 1120 985
rect 1140 965 1160 985
rect 1180 965 1200 985
rect 1220 965 1240 985
rect 1260 965 1280 985
rect 1300 965 1320 985
rect 1340 965 1360 985
rect 1380 965 1400 985
rect 1420 965 1440 985
rect 1460 965 1470 985
rect 670 821 1470 965
rect 670 801 680 821
rect 700 801 720 821
rect 740 801 760 821
rect 780 801 800 821
rect 820 801 840 821
rect 860 801 880 821
rect 900 801 920 821
rect 940 801 960 821
rect 980 801 1000 821
rect 1020 801 1040 821
rect 1060 801 1080 821
rect 1100 801 1120 821
rect 1140 801 1160 821
rect 1180 801 1200 821
rect 1220 801 1240 821
rect 1260 801 1280 821
rect 1300 801 1320 821
rect 1340 801 1360 821
rect 1380 801 1400 821
rect 1420 801 1440 821
rect 1460 801 1470 821
rect 670 657 1470 801
rect 670 637 680 657
rect 700 637 720 657
rect 740 637 760 657
rect 780 637 800 657
rect 820 637 840 657
rect 860 637 880 657
rect 900 637 920 657
rect 940 637 960 657
rect 980 637 1000 657
rect 1020 637 1040 657
rect 1060 637 1080 657
rect 1100 637 1120 657
rect 1140 637 1160 657
rect 1180 637 1200 657
rect 1220 637 1240 657
rect 1260 637 1280 657
rect 1300 637 1320 657
rect 1340 637 1360 657
rect 1380 637 1400 657
rect 1420 637 1440 657
rect 1460 637 1470 657
rect 670 493 1470 637
rect 670 473 680 493
rect 700 473 720 493
rect 740 473 760 493
rect 780 473 800 493
rect 820 473 840 493
rect 860 473 880 493
rect 900 473 920 493
rect 940 473 960 493
rect 980 473 1000 493
rect 1020 473 1040 493
rect 1060 473 1080 493
rect 1100 473 1120 493
rect 1140 473 1160 493
rect 1180 473 1200 493
rect 1220 473 1240 493
rect 1260 473 1280 493
rect 1300 473 1320 493
rect 1340 473 1360 493
rect 1380 473 1400 493
rect 1420 473 1440 493
rect 1460 473 1470 493
rect 670 329 1470 473
rect 670 309 680 329
rect 700 309 720 329
rect 740 309 760 329
rect 780 309 800 329
rect 820 309 840 329
rect 860 309 880 329
rect 900 309 920 329
rect 940 309 960 329
rect 980 309 1000 329
rect 1020 309 1040 329
rect 1060 309 1080 329
rect 1100 309 1120 329
rect 1140 309 1160 329
rect 1180 309 1200 329
rect 1220 309 1240 329
rect 1260 309 1280 329
rect 1300 309 1320 329
rect 1340 309 1360 329
rect 1380 309 1400 329
rect 1420 309 1440 329
rect 1460 309 1470 329
rect 670 165 1470 309
rect 1750 2215 2550 2390
rect 1750 2195 1760 2215
rect 1780 2195 1800 2215
rect 1820 2195 1840 2215
rect 1860 2195 1880 2215
rect 1900 2195 1920 2215
rect 1940 2195 1960 2215
rect 1980 2195 2000 2215
rect 2020 2195 2040 2215
rect 2060 2195 2080 2215
rect 2100 2195 2120 2215
rect 2140 2195 2160 2215
rect 2180 2195 2200 2215
rect 2220 2195 2240 2215
rect 2260 2195 2280 2215
rect 2300 2195 2320 2215
rect 2340 2195 2360 2215
rect 2380 2195 2400 2215
rect 2420 2195 2440 2215
rect 2460 2195 2480 2215
rect 2500 2195 2520 2215
rect 2540 2195 2550 2215
rect 1750 2051 2550 2195
rect 1750 2031 1760 2051
rect 1780 2031 1800 2051
rect 1820 2031 1840 2051
rect 1860 2031 1880 2051
rect 1900 2031 1920 2051
rect 1940 2031 1960 2051
rect 1980 2031 2000 2051
rect 2020 2031 2040 2051
rect 2060 2031 2080 2051
rect 2100 2031 2120 2051
rect 2140 2031 2160 2051
rect 2180 2031 2200 2051
rect 2220 2031 2240 2051
rect 2260 2031 2280 2051
rect 2300 2031 2320 2051
rect 2340 2031 2360 2051
rect 2380 2031 2400 2051
rect 2420 2031 2440 2051
rect 2460 2031 2480 2051
rect 2500 2031 2520 2051
rect 2540 2031 2550 2051
rect 1750 1887 2550 2031
rect 1750 1867 1760 1887
rect 1780 1867 1800 1887
rect 1820 1867 1840 1887
rect 1860 1867 1880 1887
rect 1900 1867 1920 1887
rect 1940 1867 1960 1887
rect 1980 1867 2000 1887
rect 2020 1867 2040 1887
rect 2060 1867 2080 1887
rect 2100 1867 2120 1887
rect 2140 1867 2160 1887
rect 2180 1867 2200 1887
rect 2220 1867 2240 1887
rect 2260 1867 2280 1887
rect 2300 1867 2320 1887
rect 2340 1867 2360 1887
rect 2380 1867 2400 1887
rect 2420 1867 2440 1887
rect 2460 1867 2480 1887
rect 2500 1867 2520 1887
rect 2540 1867 2550 1887
rect 1750 1723 2550 1867
rect 1750 1703 1760 1723
rect 1780 1703 1800 1723
rect 1820 1703 1840 1723
rect 1860 1703 1880 1723
rect 1900 1703 1920 1723
rect 1940 1703 1960 1723
rect 1980 1703 2000 1723
rect 2020 1703 2040 1723
rect 2060 1703 2080 1723
rect 2100 1703 2120 1723
rect 2140 1703 2160 1723
rect 2180 1703 2200 1723
rect 2220 1703 2240 1723
rect 2260 1703 2280 1723
rect 2300 1703 2320 1723
rect 2340 1703 2360 1723
rect 2380 1703 2400 1723
rect 2420 1703 2440 1723
rect 2460 1703 2480 1723
rect 2500 1703 2520 1723
rect 2540 1703 2550 1723
rect 1750 1559 2550 1703
rect 1750 1539 1760 1559
rect 1780 1539 1800 1559
rect 1820 1539 1840 1559
rect 1860 1539 1880 1559
rect 1900 1539 1920 1559
rect 1940 1539 1960 1559
rect 1980 1539 2000 1559
rect 2020 1539 2040 1559
rect 2060 1539 2080 1559
rect 2100 1539 2120 1559
rect 2140 1539 2160 1559
rect 2180 1539 2200 1559
rect 2220 1539 2240 1559
rect 2260 1539 2280 1559
rect 2300 1539 2320 1559
rect 2340 1539 2360 1559
rect 2380 1539 2400 1559
rect 2420 1539 2440 1559
rect 2460 1539 2480 1559
rect 2500 1539 2520 1559
rect 2540 1539 2550 1559
rect 1750 1395 2550 1539
rect 1750 1375 1760 1395
rect 1780 1375 1800 1395
rect 1820 1375 1840 1395
rect 1860 1375 1880 1395
rect 1900 1375 1920 1395
rect 1940 1375 1960 1395
rect 1980 1375 2000 1395
rect 2020 1375 2040 1395
rect 2060 1375 2080 1395
rect 2100 1375 2120 1395
rect 2140 1375 2160 1395
rect 2180 1375 2200 1395
rect 2220 1375 2240 1395
rect 2260 1375 2280 1395
rect 2300 1375 2320 1395
rect 2340 1375 2360 1395
rect 2380 1375 2400 1395
rect 2420 1375 2440 1395
rect 2460 1375 2480 1395
rect 2500 1375 2520 1395
rect 2540 1375 2550 1395
rect 1750 1231 2550 1375
rect 1750 1211 1760 1231
rect 1780 1211 1800 1231
rect 1820 1211 1840 1231
rect 1860 1211 1880 1231
rect 1900 1211 1920 1231
rect 1940 1211 1960 1231
rect 1980 1211 2000 1231
rect 2020 1211 2040 1231
rect 2060 1211 2080 1231
rect 2100 1211 2120 1231
rect 2140 1211 2160 1231
rect 2180 1211 2200 1231
rect 2220 1211 2240 1231
rect 2260 1211 2280 1231
rect 2300 1211 2320 1231
rect 2340 1211 2360 1231
rect 2380 1211 2400 1231
rect 2420 1211 2440 1231
rect 2460 1211 2480 1231
rect 2500 1211 2520 1231
rect 2540 1211 2550 1231
rect 1750 1067 2550 1211
rect 1750 1047 1760 1067
rect 1780 1047 1800 1067
rect 1820 1047 1840 1067
rect 1860 1047 1880 1067
rect 1900 1047 1920 1067
rect 1940 1047 1960 1067
rect 1980 1047 2000 1067
rect 2020 1047 2040 1067
rect 2060 1047 2080 1067
rect 2100 1047 2120 1067
rect 2140 1047 2160 1067
rect 2180 1047 2200 1067
rect 2220 1047 2240 1067
rect 2260 1047 2280 1067
rect 2300 1047 2320 1067
rect 2340 1047 2360 1067
rect 2380 1047 2400 1067
rect 2420 1047 2440 1067
rect 2460 1047 2480 1067
rect 2500 1047 2520 1067
rect 2540 1047 2550 1067
rect 1750 903 2550 1047
rect 1750 883 1760 903
rect 1780 883 1800 903
rect 1820 883 1840 903
rect 1860 883 1880 903
rect 1900 883 1920 903
rect 1940 883 1960 903
rect 1980 883 2000 903
rect 2020 883 2040 903
rect 2060 883 2080 903
rect 2100 883 2120 903
rect 2140 883 2160 903
rect 2180 883 2200 903
rect 2220 883 2240 903
rect 2260 883 2280 903
rect 2300 883 2320 903
rect 2340 883 2360 903
rect 2380 883 2400 903
rect 2420 883 2440 903
rect 2460 883 2480 903
rect 2500 883 2520 903
rect 2540 883 2550 903
rect 1750 739 2550 883
rect 1750 719 1760 739
rect 1780 719 1800 739
rect 1820 719 1840 739
rect 1860 719 1880 739
rect 1900 719 1920 739
rect 1940 719 1960 739
rect 1980 719 2000 739
rect 2020 719 2040 739
rect 2060 719 2080 739
rect 2100 719 2120 739
rect 2140 719 2160 739
rect 2180 719 2200 739
rect 2220 719 2240 739
rect 2260 719 2280 739
rect 2300 719 2320 739
rect 2340 719 2360 739
rect 2380 719 2400 739
rect 2420 719 2440 739
rect 2460 719 2480 739
rect 2500 719 2520 739
rect 2540 719 2550 739
rect 1750 575 2550 719
rect 1750 555 1760 575
rect 1780 555 1800 575
rect 1820 555 1840 575
rect 1860 555 1880 575
rect 1900 555 1920 575
rect 1940 555 1960 575
rect 1980 555 2000 575
rect 2020 555 2040 575
rect 2060 555 2080 575
rect 2100 555 2120 575
rect 2140 555 2160 575
rect 2180 555 2200 575
rect 2220 555 2240 575
rect 2260 555 2280 575
rect 2300 555 2320 575
rect 2340 555 2360 575
rect 2380 555 2400 575
rect 2420 555 2440 575
rect 2460 555 2480 575
rect 2500 555 2520 575
rect 2540 555 2550 575
rect 1750 411 2550 555
rect 1750 391 1760 411
rect 1780 391 1800 411
rect 1820 391 1840 411
rect 1860 391 1880 411
rect 1900 391 1920 411
rect 1940 391 1960 411
rect 1980 391 2000 411
rect 2020 391 2040 411
rect 2060 391 2080 411
rect 2100 391 2120 411
rect 2140 391 2160 411
rect 2180 391 2200 411
rect 2220 391 2240 411
rect 2260 391 2280 411
rect 2300 391 2320 411
rect 2340 391 2360 411
rect 2380 391 2400 411
rect 2420 391 2440 411
rect 2460 391 2480 411
rect 2500 391 2520 411
rect 2540 391 2550 411
rect 1750 247 2550 391
rect 1750 227 1760 247
rect 1780 227 1800 247
rect 1820 227 1840 247
rect 1860 227 1880 247
rect 1900 227 1920 247
rect 1940 227 1960 247
rect 1980 227 2000 247
rect 2020 227 2040 247
rect 2060 227 2080 247
rect 2100 227 2120 247
rect 2140 227 2160 247
rect 2180 227 2200 247
rect 2220 227 2240 247
rect 2260 227 2280 247
rect 2300 227 2320 247
rect 2340 227 2360 247
rect 2380 227 2400 247
rect 2420 227 2440 247
rect 2460 227 2480 247
rect 2500 227 2520 247
rect 2540 227 2550 247
rect 1750 217 2550 227
rect 670 145 680 165
rect 700 145 720 165
rect 740 145 760 165
rect 780 145 800 165
rect 820 145 840 165
rect 860 145 880 165
rect 900 145 920 165
rect 940 145 960 165
rect 980 145 1000 165
rect 1020 145 1040 165
rect 1060 145 1080 165
rect 1100 145 1120 165
rect 1140 145 1160 165
rect 1180 145 1200 165
rect 1220 145 1240 165
rect 1260 145 1280 165
rect 1300 145 1320 165
rect 1340 145 1360 165
rect 1380 145 1400 165
rect 1420 145 1440 165
rect 1460 145 1470 165
rect -70 -95 85 -85
rect -70 -120 -60 -95
rect -40 -120 -20 -95
rect 0 -120 20 -95
rect 40 -120 60 -95
rect 80 -120 85 -95
rect -70 -190 85 -120
rect -70 -215 -60 -190
rect -40 -215 -20 -190
rect 0 -215 20 -190
rect 40 -215 60 -190
rect 80 -215 85 -190
rect -70 -285 85 -215
rect -70 -310 -60 -285
rect -40 -310 -20 -285
rect 0 -310 20 -285
rect 40 -310 60 -285
rect 80 -310 85 -285
rect -70 -380 85 -310
rect -70 -405 -60 -380
rect -40 -405 -20 -380
rect 0 -405 20 -380
rect 40 -405 60 -380
rect 80 -405 85 -380
rect -70 -475 85 -405
rect -70 -500 -60 -475
rect -40 -500 -20 -475
rect 0 -500 20 -475
rect 40 -500 60 -475
rect 80 -500 85 -475
rect -70 -570 85 -500
rect -70 -595 -60 -570
rect -40 -595 -20 -570
rect 0 -595 20 -570
rect 40 -595 60 -570
rect 80 -595 85 -570
rect -70 -665 85 -595
rect -70 -690 -60 -665
rect -40 -690 -20 -665
rect 0 -690 20 -665
rect 40 -690 60 -665
rect 80 -690 85 -665
rect -70 -760 85 -690
rect -70 -785 -60 -760
rect -40 -785 -20 -760
rect 0 -785 20 -760
rect 40 -785 60 -760
rect 80 -785 85 -760
rect -70 -855 85 -785
rect -70 -880 -60 -855
rect -40 -880 -20 -855
rect 0 -880 20 -855
rect 40 -880 60 -855
rect 80 -880 85 -855
rect -70 -950 85 -880
rect -70 -975 -60 -950
rect -40 -975 -20 -950
rect 0 -975 20 -950
rect 40 -975 60 -950
rect 80 -975 85 -950
rect -70 -1045 85 -975
rect -70 -1070 -60 -1045
rect -40 -1070 -20 -1045
rect 0 -1070 20 -1045
rect 40 -1070 60 -1045
rect 80 -1070 85 -1045
rect -70 -1140 85 -1070
rect -70 -1165 -60 -1140
rect -40 -1165 -20 -1140
rect 0 -1165 20 -1140
rect 40 -1165 60 -1140
rect 80 -1165 85 -1140
rect -70 -1235 85 -1165
rect -70 -1260 -60 -1235
rect -40 -1260 -20 -1235
rect 0 -1260 20 -1235
rect 40 -1260 60 -1235
rect 80 -1260 85 -1235
rect -70 -1330 85 -1260
rect -70 -1355 -60 -1330
rect -40 -1355 -20 -1330
rect 0 -1355 20 -1330
rect 40 -1355 60 -1330
rect 80 -1355 85 -1330
rect -70 -1425 85 -1355
rect -70 -1450 -60 -1425
rect -40 -1450 -20 -1425
rect 0 -1450 20 -1425
rect 40 -1450 60 -1425
rect 80 -1450 85 -1425
rect -70 -1520 85 -1450
rect -70 -1545 -60 -1520
rect -40 -1545 -20 -1520
rect 0 -1545 20 -1520
rect 40 -1545 60 -1520
rect 80 -1545 85 -1520
rect -70 -1615 85 -1545
rect -70 -1640 -60 -1615
rect -40 -1640 -20 -1615
rect 0 -1640 20 -1615
rect 40 -1640 60 -1615
rect 80 -1640 85 -1615
rect -70 -1710 85 -1640
rect -70 -1735 -60 -1710
rect -40 -1735 -20 -1710
rect 0 -1735 20 -1710
rect 40 -1735 60 -1710
rect 80 -1735 85 -1710
rect -70 -1805 85 -1735
rect -70 -1830 -60 -1805
rect -40 -1830 -20 -1805
rect 0 -1830 20 -1805
rect 40 -1830 60 -1805
rect 80 -1830 85 -1805
rect -70 -1900 85 -1830
rect -70 -1925 -60 -1900
rect -40 -1925 -20 -1900
rect 0 -1925 20 -1900
rect 40 -1925 60 -1900
rect 80 -1925 85 -1900
rect -70 -1995 85 -1925
rect -70 -2020 -60 -1995
rect -40 -2020 -20 -1995
rect 0 -2020 20 -1995
rect 40 -2020 60 -1995
rect 80 -2020 85 -1995
rect -70 -2090 85 -2020
rect -70 -2115 -60 -2090
rect -40 -2115 -20 -2090
rect 0 -2115 20 -2090
rect 40 -2115 60 -2090
rect 80 -2115 85 -2090
rect -70 -2185 85 -2115
rect -70 -2210 -60 -2185
rect -40 -2210 -20 -2185
rect 0 -2210 20 -2185
rect 40 -2210 60 -2185
rect 80 -2210 85 -2185
rect -70 -2280 85 -2210
rect -70 -2305 -60 -2280
rect -40 -2305 -20 -2280
rect 0 -2305 20 -2280
rect 40 -2305 60 -2280
rect 80 -2305 85 -2280
rect -70 -2375 85 -2305
rect -70 -2400 -60 -2375
rect -40 -2400 -20 -2375
rect 0 -2400 20 -2375
rect 40 -2400 60 -2375
rect 80 -2400 85 -2375
rect -70 -2470 85 -2400
rect 670 -145 1470 145
rect 670 -165 680 -145
rect 700 -165 720 -145
rect 740 -165 760 -145
rect 780 -165 800 -145
rect 820 -165 840 -145
rect 860 -165 880 -145
rect 900 -165 920 -145
rect 940 -165 960 -145
rect 980 -165 1000 -145
rect 1020 -165 1040 -145
rect 1060 -165 1080 -145
rect 1100 -165 1120 -145
rect 1140 -165 1160 -145
rect 1180 -165 1200 -145
rect 1220 -165 1240 -145
rect 1260 -165 1280 -145
rect 1300 -165 1320 -145
rect 1340 -165 1360 -145
rect 1380 -165 1400 -145
rect 1420 -165 1440 -145
rect 1460 -165 1470 -145
rect 670 -335 1470 -165
rect 670 -355 680 -335
rect 700 -355 720 -335
rect 740 -355 760 -335
rect 780 -355 800 -335
rect 820 -355 840 -335
rect 860 -355 880 -335
rect 900 -355 920 -335
rect 940 -355 960 -335
rect 980 -355 1000 -335
rect 1020 -355 1040 -335
rect 1060 -355 1080 -335
rect 1100 -355 1120 -335
rect 1140 -355 1160 -335
rect 1180 -355 1200 -335
rect 1220 -355 1240 -335
rect 1260 -355 1280 -335
rect 1300 -355 1320 -335
rect 1340 -355 1360 -335
rect 1380 -355 1400 -335
rect 1420 -355 1440 -335
rect 1460 -355 1470 -335
rect 670 -525 1470 -355
rect 670 -545 680 -525
rect 700 -545 720 -525
rect 740 -545 760 -525
rect 780 -545 800 -525
rect 820 -545 840 -525
rect 860 -545 880 -525
rect 900 -545 920 -525
rect 940 -545 960 -525
rect 980 -545 1000 -525
rect 1020 -545 1040 -525
rect 1060 -545 1080 -525
rect 1100 -545 1120 -525
rect 1140 -545 1160 -525
rect 1180 -545 1200 -525
rect 1220 -545 1240 -525
rect 1260 -545 1280 -525
rect 1300 -545 1320 -525
rect 1340 -545 1360 -525
rect 1380 -545 1400 -525
rect 1420 -545 1440 -525
rect 1460 -545 1470 -525
rect 670 -715 1470 -545
rect 670 -735 680 -715
rect 700 -735 720 -715
rect 740 -735 760 -715
rect 780 -735 800 -715
rect 820 -735 840 -715
rect 860 -735 880 -715
rect 900 -735 920 -715
rect 940 -735 960 -715
rect 980 -735 1000 -715
rect 1020 -735 1040 -715
rect 1060 -735 1080 -715
rect 1100 -735 1120 -715
rect 1140 -735 1160 -715
rect 1180 -735 1200 -715
rect 1220 -735 1240 -715
rect 1260 -735 1280 -715
rect 1300 -735 1320 -715
rect 1340 -735 1360 -715
rect 1380 -735 1400 -715
rect 1420 -735 1440 -715
rect 1460 -735 1470 -715
rect 670 -905 1470 -735
rect 670 -925 680 -905
rect 700 -925 720 -905
rect 740 -925 760 -905
rect 780 -925 800 -905
rect 820 -925 840 -905
rect 860 -925 880 -905
rect 900 -925 920 -905
rect 940 -925 960 -905
rect 980 -925 1000 -905
rect 1020 -925 1040 -905
rect 1060 -925 1080 -905
rect 1100 -925 1120 -905
rect 1140 -925 1160 -905
rect 1180 -925 1200 -905
rect 1220 -925 1240 -905
rect 1260 -925 1280 -905
rect 1300 -925 1320 -905
rect 1340 -925 1360 -905
rect 1380 -925 1400 -905
rect 1420 -925 1440 -905
rect 1460 -925 1470 -905
rect 670 -1095 1470 -925
rect 670 -1115 680 -1095
rect 700 -1115 720 -1095
rect 740 -1115 760 -1095
rect 780 -1115 800 -1095
rect 820 -1115 840 -1095
rect 860 -1115 880 -1095
rect 900 -1115 920 -1095
rect 940 -1115 960 -1095
rect 980 -1115 1000 -1095
rect 1020 -1115 1040 -1095
rect 1060 -1115 1080 -1095
rect 1100 -1115 1120 -1095
rect 1140 -1115 1160 -1095
rect 1180 -1115 1200 -1095
rect 1220 -1115 1240 -1095
rect 1260 -1115 1280 -1095
rect 1300 -1115 1320 -1095
rect 1340 -1115 1360 -1095
rect 1380 -1115 1400 -1095
rect 1420 -1115 1440 -1095
rect 1460 -1115 1470 -1095
rect 670 -1285 1470 -1115
rect 670 -1305 680 -1285
rect 700 -1305 720 -1285
rect 740 -1305 760 -1285
rect 780 -1305 800 -1285
rect 820 -1305 840 -1285
rect 860 -1305 880 -1285
rect 900 -1305 920 -1285
rect 940 -1305 960 -1285
rect 980 -1305 1000 -1285
rect 1020 -1305 1040 -1285
rect 1060 -1305 1080 -1285
rect 1100 -1305 1120 -1285
rect 1140 -1305 1160 -1285
rect 1180 -1305 1200 -1285
rect 1220 -1305 1240 -1285
rect 1260 -1305 1280 -1285
rect 1300 -1305 1320 -1285
rect 1340 -1305 1360 -1285
rect 1380 -1305 1400 -1285
rect 1420 -1305 1440 -1285
rect 1460 -1305 1470 -1285
rect 670 -1475 1470 -1305
rect 670 -1495 680 -1475
rect 700 -1495 720 -1475
rect 740 -1495 760 -1475
rect 780 -1495 800 -1475
rect 820 -1495 840 -1475
rect 860 -1495 880 -1475
rect 900 -1495 920 -1475
rect 940 -1495 960 -1475
rect 980 -1495 1000 -1475
rect 1020 -1495 1040 -1475
rect 1060 -1495 1080 -1475
rect 1100 -1495 1120 -1475
rect 1140 -1495 1160 -1475
rect 1180 -1495 1200 -1475
rect 1220 -1495 1240 -1475
rect 1260 -1495 1280 -1475
rect 1300 -1495 1320 -1475
rect 1340 -1495 1360 -1475
rect 1380 -1495 1400 -1475
rect 1420 -1495 1440 -1475
rect 1460 -1495 1470 -1475
rect 670 -1665 1470 -1495
rect 670 -1685 680 -1665
rect 700 -1685 720 -1665
rect 740 -1685 760 -1665
rect 780 -1685 800 -1665
rect 820 -1685 840 -1665
rect 860 -1685 880 -1665
rect 900 -1685 920 -1665
rect 940 -1685 960 -1665
rect 980 -1685 1000 -1665
rect 1020 -1685 1040 -1665
rect 1060 -1685 1080 -1665
rect 1100 -1685 1120 -1665
rect 1140 -1685 1160 -1665
rect 1180 -1685 1200 -1665
rect 1220 -1685 1240 -1665
rect 1260 -1685 1280 -1665
rect 1300 -1685 1320 -1665
rect 1340 -1685 1360 -1665
rect 1380 -1685 1400 -1665
rect 1420 -1685 1440 -1665
rect 1460 -1685 1470 -1665
rect 670 -1855 1470 -1685
rect 670 -1875 680 -1855
rect 700 -1875 720 -1855
rect 740 -1875 760 -1855
rect 780 -1875 800 -1855
rect 820 -1875 840 -1855
rect 860 -1875 880 -1855
rect 900 -1875 920 -1855
rect 940 -1875 960 -1855
rect 980 -1875 1000 -1855
rect 1020 -1875 1040 -1855
rect 1060 -1875 1080 -1855
rect 1100 -1875 1120 -1855
rect 1140 -1875 1160 -1855
rect 1180 -1875 1200 -1855
rect 1220 -1875 1240 -1855
rect 1260 -1875 1280 -1855
rect 1300 -1875 1320 -1855
rect 1340 -1875 1360 -1855
rect 1380 -1875 1400 -1855
rect 1420 -1875 1440 -1855
rect 1460 -1875 1470 -1855
rect 670 -2045 1470 -1875
rect 670 -2065 680 -2045
rect 700 -2065 720 -2045
rect 740 -2065 760 -2045
rect 780 -2065 800 -2045
rect 820 -2065 840 -2045
rect 860 -2065 880 -2045
rect 900 -2065 920 -2045
rect 940 -2065 960 -2045
rect 980 -2065 1000 -2045
rect 1020 -2065 1040 -2045
rect 1060 -2065 1080 -2045
rect 1100 -2065 1120 -2045
rect 1140 -2065 1160 -2045
rect 1180 -2065 1200 -2045
rect 1220 -2065 1240 -2045
rect 1260 -2065 1280 -2045
rect 1300 -2065 1320 -2045
rect 1340 -2065 1360 -2045
rect 1380 -2065 1400 -2045
rect 1420 -2065 1440 -2045
rect 1460 -2065 1470 -2045
rect 670 -2235 1470 -2065
rect 670 -2255 680 -2235
rect 700 -2255 720 -2235
rect 740 -2255 760 -2235
rect 780 -2255 800 -2235
rect 820 -2255 840 -2235
rect 860 -2255 880 -2235
rect 900 -2255 920 -2235
rect 940 -2255 960 -2235
rect 980 -2255 1000 -2235
rect 1020 -2255 1040 -2235
rect 1060 -2255 1080 -2235
rect 1100 -2255 1120 -2235
rect 1140 -2255 1160 -2235
rect 1180 -2255 1200 -2235
rect 1220 -2255 1240 -2235
rect 1260 -2255 1280 -2235
rect 1300 -2255 1320 -2235
rect 1340 -2255 1360 -2235
rect 1380 -2255 1400 -2235
rect 1420 -2255 1440 -2235
rect 1460 -2255 1470 -2235
rect 670 -2425 1470 -2255
rect 670 -2445 680 -2425
rect 700 -2445 720 -2425
rect 740 -2445 760 -2425
rect 780 -2445 800 -2425
rect 820 -2445 840 -2425
rect 860 -2445 880 -2425
rect 900 -2445 920 -2425
rect 940 -2445 960 -2425
rect 980 -2445 1000 -2425
rect 1020 -2445 1040 -2425
rect 1060 -2445 1080 -2425
rect 1100 -2445 1120 -2425
rect 1140 -2445 1160 -2425
rect 1180 -2445 1200 -2425
rect 1220 -2445 1240 -2425
rect 1260 -2445 1280 -2425
rect 1300 -2445 1320 -2425
rect 1340 -2445 1360 -2425
rect 1380 -2445 1400 -2425
rect 1420 -2445 1440 -2425
rect 1460 -2445 1470 -2425
rect 670 -2455 1470 -2445
rect 1750 95 2675 105
rect 1750 75 1760 95
rect 1780 75 1800 95
rect 1820 75 1840 95
rect 1860 75 1880 95
rect 1900 75 1920 95
rect 1940 75 1960 95
rect 1980 75 2000 95
rect 2020 75 2040 95
rect 2060 75 2080 95
rect 2100 75 2120 95
rect 2140 75 2160 95
rect 2180 75 2200 95
rect 2220 75 2240 95
rect 2260 75 2280 95
rect 2300 75 2320 95
rect 2340 75 2360 95
rect 2380 75 2400 95
rect 2420 75 2440 95
rect 2460 75 2480 95
rect 2500 75 2520 95
rect 2540 75 2560 95
rect 2580 75 2600 95
rect 2620 75 2640 95
rect 2660 75 2675 95
rect 1750 50 2675 75
rect 1750 -10 2550 50
rect 1750 -30 1760 -10
rect 1780 -30 1800 -10
rect 1820 -30 1840 -10
rect 1860 -30 1880 -10
rect 1900 -30 1920 -10
rect 1940 -30 1960 -10
rect 1980 -30 2000 -10
rect 2020 -30 2040 -10
rect 2060 -30 2080 -10
rect 2100 -30 2120 -10
rect 2140 -30 2160 -10
rect 2180 -30 2200 -10
rect 2220 -30 2240 -10
rect 2260 -30 2280 -10
rect 2300 -30 2320 -10
rect 2340 -30 2360 -10
rect 2380 -30 2400 -10
rect 2420 -30 2440 -10
rect 2460 -30 2480 -10
rect 2500 -30 2520 -10
rect 2540 -30 2550 -10
rect 1750 -50 2550 -30
rect 1750 -70 1760 -50
rect 1780 -70 1800 -50
rect 1820 -70 1840 -50
rect 1860 -70 1880 -50
rect 1900 -70 1920 -50
rect 1940 -70 1960 -50
rect 1980 -70 2000 -50
rect 2020 -70 2040 -50
rect 2060 -70 2080 -50
rect 2100 -70 2120 -50
rect 2140 -70 2160 -50
rect 2180 -70 2200 -50
rect 2220 -70 2240 -50
rect 2260 -70 2280 -50
rect 2300 -70 2320 -50
rect 2340 -70 2360 -50
rect 2380 -70 2400 -50
rect 2420 -70 2440 -50
rect 2460 -70 2480 -50
rect 2500 -70 2520 -50
rect 2540 -70 2550 -50
rect 1750 -240 2550 -70
rect 1750 -260 1760 -240
rect 1780 -260 1800 -240
rect 1820 -260 1840 -240
rect 1860 -260 1880 -240
rect 1900 -260 1920 -240
rect 1940 -260 1960 -240
rect 1980 -260 2000 -240
rect 2020 -260 2040 -240
rect 2060 -260 2080 -240
rect 2100 -260 2120 -240
rect 2140 -260 2160 -240
rect 2180 -260 2200 -240
rect 2220 -260 2240 -240
rect 2260 -260 2280 -240
rect 2300 -260 2320 -240
rect 2340 -260 2360 -240
rect 2380 -260 2400 -240
rect 2420 -260 2440 -240
rect 2460 -260 2480 -240
rect 2500 -260 2520 -240
rect 2540 -260 2550 -240
rect 1750 -430 2550 -260
rect 1750 -450 1760 -430
rect 1780 -450 1800 -430
rect 1820 -450 1840 -430
rect 1860 -450 1880 -430
rect 1900 -450 1920 -430
rect 1940 -450 1960 -430
rect 1980 -450 2000 -430
rect 2020 -450 2040 -430
rect 2060 -450 2080 -430
rect 2100 -450 2120 -430
rect 2140 -450 2160 -430
rect 2180 -450 2200 -430
rect 2220 -450 2240 -430
rect 2260 -450 2280 -430
rect 2300 -450 2320 -430
rect 2340 -450 2360 -430
rect 2380 -450 2400 -430
rect 2420 -450 2440 -430
rect 2460 -450 2480 -430
rect 2500 -450 2520 -430
rect 2540 -450 2550 -430
rect 1750 -620 2550 -450
rect 1750 -640 1760 -620
rect 1780 -640 1800 -620
rect 1820 -640 1840 -620
rect 1860 -640 1880 -620
rect 1900 -640 1920 -620
rect 1940 -640 1960 -620
rect 1980 -640 2000 -620
rect 2020 -640 2040 -620
rect 2060 -640 2080 -620
rect 2100 -640 2120 -620
rect 2140 -640 2160 -620
rect 2180 -640 2200 -620
rect 2220 -640 2240 -620
rect 2260 -640 2280 -620
rect 2300 -640 2320 -620
rect 2340 -640 2360 -620
rect 2380 -640 2400 -620
rect 2420 -640 2440 -620
rect 2460 -640 2480 -620
rect 2500 -640 2520 -620
rect 2540 -640 2550 -620
rect 1750 -810 2550 -640
rect 1750 -830 1760 -810
rect 1780 -830 1800 -810
rect 1820 -830 1840 -810
rect 1860 -830 1880 -810
rect 1900 -830 1920 -810
rect 1940 -830 1960 -810
rect 1980 -830 2000 -810
rect 2020 -830 2040 -810
rect 2060 -830 2080 -810
rect 2100 -830 2120 -810
rect 2140 -830 2160 -810
rect 2180 -830 2200 -810
rect 2220 -830 2240 -810
rect 2260 -830 2280 -810
rect 2300 -830 2320 -810
rect 2340 -830 2360 -810
rect 2380 -830 2400 -810
rect 2420 -830 2440 -810
rect 2460 -830 2480 -810
rect 2500 -830 2520 -810
rect 2540 -830 2550 -810
rect 1750 -1000 2550 -830
rect 1750 -1020 1760 -1000
rect 1780 -1020 1800 -1000
rect 1820 -1020 1840 -1000
rect 1860 -1020 1880 -1000
rect 1900 -1020 1920 -1000
rect 1940 -1020 1960 -1000
rect 1980 -1020 2000 -1000
rect 2020 -1020 2040 -1000
rect 2060 -1020 2080 -1000
rect 2100 -1020 2120 -1000
rect 2140 -1020 2160 -1000
rect 2180 -1020 2200 -1000
rect 2220 -1020 2240 -1000
rect 2260 -1020 2280 -1000
rect 2300 -1020 2320 -1000
rect 2340 -1020 2360 -1000
rect 2380 -1020 2400 -1000
rect 2420 -1020 2440 -1000
rect 2460 -1020 2480 -1000
rect 2500 -1020 2520 -1000
rect 2540 -1020 2550 -1000
rect 1750 -1190 2550 -1020
rect 1750 -1210 1760 -1190
rect 1780 -1210 1800 -1190
rect 1820 -1210 1840 -1190
rect 1860 -1210 1880 -1190
rect 1900 -1210 1920 -1190
rect 1940 -1210 1960 -1190
rect 1980 -1210 2000 -1190
rect 2020 -1210 2040 -1190
rect 2060 -1210 2080 -1190
rect 2100 -1210 2120 -1190
rect 2140 -1210 2160 -1190
rect 2180 -1210 2200 -1190
rect 2220 -1210 2240 -1190
rect 2260 -1210 2280 -1190
rect 2300 -1210 2320 -1190
rect 2340 -1210 2360 -1190
rect 2380 -1210 2400 -1190
rect 2420 -1210 2440 -1190
rect 2460 -1210 2480 -1190
rect 2500 -1210 2520 -1190
rect 2540 -1210 2550 -1190
rect 1750 -1380 2550 -1210
rect 1750 -1400 1760 -1380
rect 1780 -1400 1800 -1380
rect 1820 -1400 1840 -1380
rect 1860 -1400 1880 -1380
rect 1900 -1400 1920 -1380
rect 1940 -1400 1960 -1380
rect 1980 -1400 2000 -1380
rect 2020 -1400 2040 -1380
rect 2060 -1400 2080 -1380
rect 2100 -1400 2120 -1380
rect 2140 -1400 2160 -1380
rect 2180 -1400 2200 -1380
rect 2220 -1400 2240 -1380
rect 2260 -1400 2280 -1380
rect 2300 -1400 2320 -1380
rect 2340 -1400 2360 -1380
rect 2380 -1400 2400 -1380
rect 2420 -1400 2440 -1380
rect 2460 -1400 2480 -1380
rect 2500 -1400 2520 -1380
rect 2540 -1400 2550 -1380
rect 1750 -1570 2550 -1400
rect 1750 -1590 1760 -1570
rect 1780 -1590 1800 -1570
rect 1820 -1590 1840 -1570
rect 1860 -1590 1880 -1570
rect 1900 -1590 1920 -1570
rect 1940 -1590 1960 -1570
rect 1980 -1590 2000 -1570
rect 2020 -1590 2040 -1570
rect 2060 -1590 2080 -1570
rect 2100 -1590 2120 -1570
rect 2140 -1590 2160 -1570
rect 2180 -1590 2200 -1570
rect 2220 -1590 2240 -1570
rect 2260 -1590 2280 -1570
rect 2300 -1590 2320 -1570
rect 2340 -1590 2360 -1570
rect 2380 -1590 2400 -1570
rect 2420 -1590 2440 -1570
rect 2460 -1590 2480 -1570
rect 2500 -1590 2520 -1570
rect 2540 -1590 2550 -1570
rect 1750 -1760 2550 -1590
rect 1750 -1780 1760 -1760
rect 1780 -1780 1800 -1760
rect 1820 -1780 1840 -1760
rect 1860 -1780 1880 -1760
rect 1900 -1780 1920 -1760
rect 1940 -1780 1960 -1760
rect 1980 -1780 2000 -1760
rect 2020 -1780 2040 -1760
rect 2060 -1780 2080 -1760
rect 2100 -1780 2120 -1760
rect 2140 -1780 2160 -1760
rect 2180 -1780 2200 -1760
rect 2220 -1780 2240 -1760
rect 2260 -1780 2280 -1760
rect 2300 -1780 2320 -1760
rect 2340 -1780 2360 -1760
rect 2380 -1780 2400 -1760
rect 2420 -1780 2440 -1760
rect 2460 -1780 2480 -1760
rect 2500 -1780 2520 -1760
rect 2540 -1780 2550 -1760
rect 1750 -1950 2550 -1780
rect 1750 -1970 1760 -1950
rect 1780 -1970 1800 -1950
rect 1820 -1970 1840 -1950
rect 1860 -1970 1880 -1950
rect 1900 -1970 1920 -1950
rect 1940 -1970 1960 -1950
rect 1980 -1970 2000 -1950
rect 2020 -1970 2040 -1950
rect 2060 -1970 2080 -1950
rect 2100 -1970 2120 -1950
rect 2140 -1970 2160 -1950
rect 2180 -1970 2200 -1950
rect 2220 -1970 2240 -1950
rect 2260 -1970 2280 -1950
rect 2300 -1970 2320 -1950
rect 2340 -1970 2360 -1950
rect 2380 -1970 2400 -1950
rect 2420 -1970 2440 -1950
rect 2460 -1970 2480 -1950
rect 2500 -1970 2520 -1950
rect 2540 -1970 2550 -1950
rect 1750 -2140 2550 -1970
rect 1750 -2160 1760 -2140
rect 1780 -2160 1800 -2140
rect 1820 -2160 1840 -2140
rect 1860 -2160 1880 -2140
rect 1900 -2160 1920 -2140
rect 1940 -2160 1960 -2140
rect 1980 -2160 2000 -2140
rect 2020 -2160 2040 -2140
rect 2060 -2160 2080 -2140
rect 2100 -2160 2120 -2140
rect 2140 -2160 2160 -2140
rect 2180 -2160 2200 -2140
rect 2220 -2160 2240 -2140
rect 2260 -2160 2280 -2140
rect 2300 -2160 2320 -2140
rect 2340 -2160 2360 -2140
rect 2380 -2160 2400 -2140
rect 2420 -2160 2440 -2140
rect 2460 -2160 2480 -2140
rect 2500 -2160 2520 -2140
rect 2540 -2160 2550 -2140
rect 1750 -2330 2550 -2160
rect 1750 -2350 1760 -2330
rect 1780 -2350 1800 -2330
rect 1820 -2350 1840 -2330
rect 1860 -2350 1880 -2330
rect 1900 -2350 1920 -2330
rect 1940 -2350 1960 -2330
rect 1980 -2350 2000 -2330
rect 2020 -2350 2040 -2330
rect 2060 -2350 2080 -2330
rect 2100 -2350 2120 -2330
rect 2140 -2350 2160 -2330
rect 2180 -2350 2200 -2330
rect 2220 -2350 2240 -2330
rect 2260 -2350 2280 -2330
rect 2300 -2350 2320 -2330
rect 2340 -2350 2360 -2330
rect 2380 -2350 2400 -2330
rect 2420 -2350 2440 -2330
rect 2460 -2350 2480 -2330
rect 2500 -2350 2520 -2330
rect 2540 -2350 2550 -2330
rect -70 -2495 -60 -2470
rect -40 -2495 -20 -2470
rect 0 -2495 20 -2470
rect 40 -2495 60 -2470
rect 80 -2495 85 -2470
rect -70 -2505 85 -2495
rect 1750 -2520 2550 -2350
rect 1750 -2540 1760 -2520
rect 1780 -2540 1800 -2520
rect 1820 -2540 1840 -2520
rect 1860 -2540 1880 -2520
rect 1900 -2540 1920 -2520
rect 1940 -2540 1960 -2520
rect 1980 -2540 2000 -2520
rect 2020 -2540 2040 -2520
rect 2060 -2540 2080 -2520
rect 2100 -2540 2120 -2520
rect 2140 -2540 2160 -2520
rect 2180 -2540 2200 -2520
rect 2220 -2540 2240 -2520
rect 2260 -2540 2280 -2520
rect 2300 -2540 2320 -2520
rect 2340 -2540 2360 -2520
rect 2380 -2540 2400 -2520
rect 2420 -2540 2440 -2520
rect 2460 -2540 2480 -2520
rect 2500 -2540 2520 -2520
rect 2540 -2540 2550 -2520
rect 1750 -2560 2550 -2540
rect 1750 -2580 1760 -2560
rect 1780 -2580 1800 -2560
rect 1820 -2580 1840 -2560
rect 1860 -2580 1880 -2560
rect 1900 -2580 1920 -2560
rect 1940 -2580 1960 -2560
rect 1980 -2580 2000 -2560
rect 2020 -2580 2040 -2560
rect 2060 -2580 2080 -2560
rect 2100 -2580 2120 -2560
rect 2140 -2580 2160 -2560
rect 2180 -2580 2200 -2560
rect 2220 -2580 2240 -2560
rect 2260 -2580 2280 -2560
rect 2300 -2580 2320 -2560
rect 2340 -2580 2360 -2560
rect 2380 -2580 2400 -2560
rect 2420 -2580 2440 -2560
rect 2460 -2580 2480 -2560
rect 2500 -2580 2520 -2560
rect 2540 -2580 2550 -2560
rect 1750 -2630 2550 -2580
<< labels >>
rlabel metal1 9 1164 9 1164 1 g_u
port 3 n
rlabel metal1 -59 -1294 -59 -1294 1 g_d
port 4 n
rlabel metal1 1070 20 1070 20 1 Vout
port 1 n
rlabel metal1 2170 -2610 2170 -2610 1 GND
port 8 n
rlabel metal1 2160 2385 2160 2385 1 VDD
port 9 n
<< end >>
