magic
tech sky130A
timestamp 1634684585
<< nwell >>
rect -565 1990 -560 2035
rect -565 1930 -560 1970
rect -565 1860 -560 1900
rect -565 1795 -560 1840
rect -240 1795 -235 2035
<< poly >>
rect -565 2025 -235 2035
rect -565 2005 -555 2025
rect -530 2005 -510 2025
rect -490 2005 -470 2025
rect -450 2005 -430 2025
rect -410 2005 -390 2025
rect -370 2005 -350 2025
rect -330 2005 -310 2025
rect -290 2005 -270 2025
rect -245 2005 -235 2025
rect -565 1995 -235 2005
rect -565 1960 -235 1970
rect -565 1940 -555 1960
rect -530 1940 -510 1960
rect -490 1940 -470 1960
rect -450 1940 -430 1960
rect -410 1940 -390 1960
rect -370 1940 -350 1960
rect -330 1940 -310 1960
rect -290 1940 -270 1960
rect -245 1940 -235 1960
rect -565 1930 -235 1940
rect -565 1890 -235 1900
rect -565 1870 -555 1890
rect -530 1870 -510 1890
rect -490 1870 -470 1890
rect -450 1870 -430 1890
rect -410 1870 -390 1890
rect -370 1870 -350 1890
rect -330 1870 -310 1890
rect -290 1870 -270 1890
rect -245 1870 -235 1890
rect -565 1860 -235 1870
rect -565 1825 -235 1835
rect -565 1805 -555 1825
rect -530 1805 -510 1825
rect -490 1805 -470 1825
rect -450 1805 -430 1825
rect -410 1805 -390 1825
rect -370 1805 -350 1825
rect -330 1805 -310 1825
rect -290 1805 -270 1825
rect -245 1805 -235 1825
rect -565 1795 -235 1805
<< polycont >>
rect -555 2005 -530 2025
rect -510 2005 -490 2025
rect -470 2005 -450 2025
rect -430 2005 -410 2025
rect -390 2005 -370 2025
rect -350 2005 -330 2025
rect -310 2005 -290 2025
rect -270 2005 -245 2025
rect -555 1940 -530 1960
rect -510 1940 -490 1960
rect -470 1940 -450 1960
rect -430 1940 -410 1960
rect -390 1940 -370 1960
rect -350 1940 -330 1960
rect -310 1940 -290 1960
rect -270 1940 -245 1960
rect -555 1870 -530 1890
rect -510 1870 -490 1890
rect -470 1870 -450 1890
rect -430 1870 -410 1890
rect -390 1870 -370 1890
rect -350 1870 -330 1890
rect -310 1870 -290 1890
rect -270 1870 -245 1890
rect -555 1805 -530 1825
rect -510 1805 -490 1825
rect -470 1805 -450 1825
rect -430 1805 -410 1825
rect -390 1805 -370 1825
rect -350 1805 -330 1825
rect -310 1805 -290 1825
rect -270 1805 -245 1825
<< xpolycontact >>
rect -710 630 -470 771
rect -329 630 -90 771
<< xpolyres >>
rect -470 630 -329 771
<< locali >>
rect -555 2025 -245 2035
rect -530 2005 -510 2025
rect -490 2005 -470 2025
rect -450 2005 -430 2025
rect -410 2005 -390 2025
rect -370 2005 -350 2025
rect -330 2005 -310 2025
rect -290 2005 -270 2025
rect -555 1995 -245 2005
rect -555 1960 -245 1970
rect -530 1940 -510 1960
rect -490 1940 -470 1960
rect -450 1940 -430 1960
rect -410 1940 -390 1960
rect -370 1940 -350 1960
rect -330 1940 -310 1960
rect -290 1940 -270 1960
rect -555 1930 -245 1940
rect -555 1890 -245 1900
rect -530 1870 -510 1890
rect -490 1870 -470 1890
rect -450 1870 -430 1890
rect -410 1870 -390 1890
rect -370 1870 -350 1890
rect -330 1870 -310 1890
rect -290 1870 -270 1890
rect -555 1860 -245 1870
rect -555 1825 -245 1835
rect -530 1805 -510 1825
rect -490 1805 -470 1825
rect -450 1805 -430 1825
rect -410 1805 -390 1825
rect -370 1805 -350 1825
rect -330 1805 -310 1825
rect -290 1805 -270 1825
rect -555 1795 -245 1805
<< viali >>
rect -550 2005 -530 2025
rect -510 2005 -490 2025
rect -470 2005 -450 2025
rect -430 2005 -410 2025
rect -390 2005 -370 2025
rect -350 2005 -330 2025
rect -310 2005 -290 2025
rect -270 2005 -250 2025
rect -550 1940 -530 1960
rect -510 1940 -490 1960
rect -470 1940 -450 1960
rect -430 1940 -410 1960
rect -390 1940 -370 1960
rect -350 1940 -330 1960
rect -310 1940 -290 1960
rect -270 1940 -250 1960
rect -550 1870 -530 1890
rect -510 1870 -490 1890
rect -470 1870 -450 1890
rect -430 1870 -410 1890
rect -390 1870 -370 1890
rect -350 1870 -330 1890
rect -310 1870 -290 1890
rect -270 1870 -250 1890
rect -550 1805 -530 1825
rect -510 1805 -490 1825
rect -470 1805 -450 1825
rect -430 1805 -410 1825
rect -390 1805 -370 1825
rect -350 1805 -330 1825
rect -310 1805 -290 1825
rect -270 1805 -250 1825
rect -700 730 -680 750
rect -660 730 -640 750
rect -620 730 -600 750
rect -580 730 -560 750
rect -540 730 -520 750
rect -500 730 -480 750
rect -700 690 -680 710
rect -660 690 -640 710
rect -620 690 -600 710
rect -580 690 -560 710
rect -540 690 -520 710
rect -500 690 -480 710
rect -700 650 -680 670
rect -660 650 -640 670
rect -620 650 -600 670
rect -580 650 -560 670
rect -540 650 -520 670
rect -500 650 -480 670
rect -320 730 -300 750
rect -280 730 -260 750
rect -240 730 -220 750
rect -200 730 -180 750
rect -160 730 -140 750
rect -120 730 -100 750
rect -320 690 -300 710
rect -280 690 -260 710
rect -240 690 -220 710
rect -200 690 -180 710
rect -160 690 -140 710
rect -120 690 -100 710
rect -320 650 -300 670
rect -280 650 -260 670
rect -240 650 -220 670
rect -200 650 -180 670
rect -160 650 -140 670
rect -120 650 -100 670
<< metal1 >>
rect -1010 2120 -1000 2130
rect 200 2120 210 2130
rect -565 2025 -235 2035
rect -565 2005 -550 2025
rect -530 2005 -510 2025
rect -490 2005 -470 2025
rect -450 2005 -430 2025
rect -410 2005 -390 2025
rect -370 2005 -350 2025
rect -330 2005 -310 2025
rect -290 2005 -270 2025
rect -250 2005 -235 2025
rect -565 1960 -235 2005
rect -565 1940 -550 1960
rect -530 1940 -510 1960
rect -490 1940 -470 1960
rect -450 1940 -430 1960
rect -410 1940 -390 1960
rect -370 1940 -350 1960
rect -330 1940 -310 1960
rect -290 1940 -270 1960
rect -250 1940 -235 1960
rect -565 1890 -235 1940
rect -565 1870 -550 1890
rect -530 1870 -510 1890
rect -490 1870 -470 1890
rect -450 1870 -430 1890
rect -410 1870 -390 1890
rect -370 1870 -350 1890
rect -330 1870 -310 1890
rect -290 1870 -270 1890
rect -250 1870 -235 1890
rect -565 1825 -235 1870
rect -565 1805 -550 1825
rect -530 1805 -510 1825
rect -490 1805 -470 1825
rect -450 1805 -430 1825
rect -410 1805 -390 1825
rect -370 1805 -350 1825
rect -330 1805 -310 1825
rect -290 1805 -270 1825
rect -250 1805 -235 1825
rect -565 1795 -235 1805
rect -310 1740 -235 1795
rect -1375 1710 -1365 1720
rect -310 1715 450 1740
rect -1955 1115 -1945 1125
rect 1145 1120 1155 1130
rect -950 750 -470 771
rect -950 730 -700 750
rect -680 730 -660 750
rect -640 730 -620 750
rect -600 730 -580 750
rect -560 730 -540 750
rect -520 730 -500 750
rect -480 730 -470 750
rect -950 710 -470 730
rect -950 690 -700 710
rect -680 690 -660 710
rect -640 690 -620 710
rect -600 690 -580 710
rect -560 690 -540 710
rect -520 690 -500 710
rect -480 690 -470 710
rect -950 670 -470 690
rect -950 650 -700 670
rect -680 650 -660 670
rect -640 650 -620 670
rect -600 650 -580 670
rect -560 650 -540 670
rect -520 650 -500 670
rect -480 650 -470 670
rect -950 630 -470 650
rect -329 750 125 771
rect -329 730 -320 750
rect -300 730 -280 750
rect -260 730 -240 750
rect -220 730 -200 750
rect -180 730 -160 750
rect -140 730 -120 750
rect -100 730 125 750
rect -329 710 125 730
rect -329 690 -320 710
rect -300 690 -280 710
rect -260 690 -240 710
rect -220 690 -200 710
rect -180 690 -160 710
rect -140 690 -120 710
rect -100 690 125 710
rect -329 670 125 690
rect -329 650 -320 670
rect -300 650 -280 670
rect -260 650 -240 670
rect -220 650 -200 670
rect -180 650 -160 670
rect -140 650 -120 670
rect -100 650 125 670
rect -329 630 125 650
rect -500 45 -300 495
rect -1535 -15 -1525 -5
rect 705 -15 715 -5
use cmfb_half  cmfb_half_0
timestamp 1634684585
transform 1 0 -35 0 1 1205
box -310 -1220 1190 930
use cmfb_half  cmfb_half_1
timestamp 1634684585
transform -1 0 -765 0 1 1205
box -310 -1220 1190 930
<< labels >>
rlabel metal1 -405 275 -405 275 1 Vb3
port 13 n
rlabel metal1 -1950 1120 -1950 1120 1 Vref
port 14 n
rlabel metal1 1150 1125 1150 1125 1 Vcm
port 15 n
rlabel metal1 710 -10 710 -10 1 GND#1
port 16 n
rlabel metal1 -1530 -10 -1530 -10 1 GND
port 17 n
rlabel metal1 -1005 2125 -1005 2125 1 VDD
port 18 n
rlabel metal1 -1370 1715 -1370 1715 1 Vcmfb
port 20 n
rlabel metal1 205 2125 205 2125 1 VDD
port 18 n
<< end >>
