magic
tech sky130A
timestamp 1634684585
<< nwell >>
rect -205 530 885 930
<< nmos >>
rect 15 430 1015 450
rect 15 360 1015 380
rect 15 290 1015 310
rect 15 220 1015 240
rect 15 150 1015 170
rect 15 80 1015 100
rect 15 10 1015 30
rect 15 -60 1015 -40
rect 15 -130 1015 -110
rect 15 -200 1015 -180
rect 15 -270 1015 -250
rect 15 -340 1015 -320
rect 15 -410 1015 -390
rect 15 -480 1015 -460
rect 15 -550 1015 -530
rect -135 -760 1165 -710
rect -135 -860 1165 -810
rect -135 -960 1165 -910
rect -135 -1060 1165 -1010
rect -135 -1160 1165 -1110
<< pmos >>
rect -185 805 865 825
rect -185 735 865 755
rect -185 665 865 685
rect -185 595 865 615
<< ndiff >>
rect 15 485 1015 495
rect 15 465 30 485
rect 65 465 85 485
rect 105 465 125 485
rect 145 465 165 485
rect 185 465 205 485
rect 225 465 245 485
rect 265 465 285 485
rect 305 465 325 485
rect 345 465 365 485
rect 385 465 405 485
rect 425 465 445 485
rect 465 465 485 485
rect 505 465 525 485
rect 545 465 565 485
rect 585 465 605 485
rect 625 465 645 485
rect 665 465 685 485
rect 705 465 725 485
rect 745 465 765 485
rect 785 465 805 485
rect 825 465 845 485
rect 865 465 885 485
rect 905 465 925 485
rect 945 465 965 485
rect 1000 465 1015 485
rect 15 450 1015 465
rect 15 415 1015 430
rect 15 395 30 415
rect 65 395 85 415
rect 105 395 125 415
rect 145 395 165 415
rect 185 395 205 415
rect 225 395 245 415
rect 265 395 285 415
rect 305 395 325 415
rect 345 395 365 415
rect 385 395 405 415
rect 425 395 445 415
rect 465 395 485 415
rect 505 395 525 415
rect 545 395 565 415
rect 585 395 605 415
rect 625 395 645 415
rect 665 395 685 415
rect 705 395 725 415
rect 745 395 765 415
rect 785 395 805 415
rect 825 395 845 415
rect 865 395 885 415
rect 905 395 925 415
rect 945 395 965 415
rect 1000 395 1015 415
rect 15 380 1015 395
rect 15 345 1015 360
rect 15 325 30 345
rect 65 325 85 345
rect 105 325 125 345
rect 145 325 165 345
rect 185 325 205 345
rect 225 325 245 345
rect 265 325 285 345
rect 305 325 325 345
rect 345 325 365 345
rect 385 325 405 345
rect 425 325 445 345
rect 465 325 485 345
rect 505 325 525 345
rect 545 325 565 345
rect 585 325 605 345
rect 625 325 645 345
rect 665 325 685 345
rect 705 325 725 345
rect 745 325 765 345
rect 785 325 805 345
rect 825 325 845 345
rect 865 325 885 345
rect 905 325 925 345
rect 945 325 965 345
rect 1000 325 1015 345
rect 15 310 1015 325
rect 15 275 1015 290
rect 15 255 30 275
rect 65 255 85 275
rect 105 255 125 275
rect 145 255 165 275
rect 185 255 205 275
rect 225 255 245 275
rect 265 255 285 275
rect 305 255 325 275
rect 345 255 365 275
rect 385 255 405 275
rect 425 255 445 275
rect 465 255 485 275
rect 505 255 525 275
rect 545 255 565 275
rect 585 255 605 275
rect 625 255 645 275
rect 665 255 685 275
rect 705 255 725 275
rect 745 255 765 275
rect 785 255 805 275
rect 825 255 845 275
rect 865 255 885 275
rect 905 255 925 275
rect 945 255 965 275
rect 1000 255 1015 275
rect 15 240 1015 255
rect 15 205 1015 220
rect 15 185 30 205
rect 65 185 85 205
rect 105 185 125 205
rect 145 185 165 205
rect 185 185 205 205
rect 225 185 245 205
rect 265 185 285 205
rect 305 185 325 205
rect 345 185 365 205
rect 385 185 405 205
rect 425 185 445 205
rect 465 185 485 205
rect 505 185 525 205
rect 545 185 565 205
rect 585 185 605 205
rect 625 185 645 205
rect 665 185 685 205
rect 705 185 725 205
rect 745 185 765 205
rect 785 185 805 205
rect 825 185 845 205
rect 865 185 885 205
rect 905 185 925 205
rect 945 185 965 205
rect 1000 185 1015 205
rect 15 170 1015 185
rect 15 135 1015 150
rect 15 115 30 135
rect 65 115 85 135
rect 105 115 125 135
rect 145 115 165 135
rect 185 115 205 135
rect 225 115 245 135
rect 265 115 285 135
rect 305 115 325 135
rect 345 115 365 135
rect 385 115 405 135
rect 425 115 445 135
rect 465 115 485 135
rect 505 115 525 135
rect 545 115 565 135
rect 585 115 605 135
rect 625 115 645 135
rect 665 115 685 135
rect 705 115 725 135
rect 745 115 765 135
rect 785 115 805 135
rect 825 115 845 135
rect 865 115 885 135
rect 905 115 925 135
rect 945 115 965 135
rect 1000 115 1015 135
rect 15 100 1015 115
rect 15 65 1015 80
rect 15 45 30 65
rect 65 45 85 65
rect 105 45 125 65
rect 145 45 165 65
rect 185 45 205 65
rect 225 45 245 65
rect 265 45 285 65
rect 305 45 325 65
rect 345 45 365 65
rect 385 45 405 65
rect 425 45 445 65
rect 465 45 485 65
rect 505 45 525 65
rect 545 45 565 65
rect 585 45 605 65
rect 625 45 645 65
rect 665 45 685 65
rect 705 45 725 65
rect 745 45 765 65
rect 785 45 805 65
rect 825 45 845 65
rect 865 45 885 65
rect 905 45 925 65
rect 945 45 965 65
rect 1000 45 1015 65
rect 15 30 1015 45
rect 15 -5 1015 10
rect 15 -25 30 -5
rect 65 -25 85 -5
rect 105 -25 125 -5
rect 145 -25 165 -5
rect 185 -25 205 -5
rect 225 -25 245 -5
rect 265 -25 285 -5
rect 305 -25 325 -5
rect 345 -25 365 -5
rect 385 -25 405 -5
rect 425 -25 445 -5
rect 465 -25 485 -5
rect 505 -25 525 -5
rect 545 -25 565 -5
rect 585 -25 605 -5
rect 625 -25 645 -5
rect 665 -25 685 -5
rect 705 -25 725 -5
rect 745 -25 765 -5
rect 785 -25 805 -5
rect 825 -25 845 -5
rect 865 -25 885 -5
rect 905 -25 925 -5
rect 945 -25 965 -5
rect 1000 -25 1015 -5
rect 15 -40 1015 -25
rect 15 -75 1015 -60
rect 15 -95 30 -75
rect 65 -95 85 -75
rect 105 -95 125 -75
rect 145 -95 165 -75
rect 185 -95 205 -75
rect 225 -95 245 -75
rect 265 -95 285 -75
rect 305 -95 325 -75
rect 345 -95 365 -75
rect 385 -95 405 -75
rect 425 -95 445 -75
rect 465 -95 485 -75
rect 505 -95 525 -75
rect 545 -95 565 -75
rect 585 -95 605 -75
rect 625 -95 645 -75
rect 665 -95 685 -75
rect 705 -95 725 -75
rect 745 -95 765 -75
rect 785 -95 805 -75
rect 825 -95 845 -75
rect 865 -95 885 -75
rect 905 -95 925 -75
rect 945 -95 965 -75
rect 1000 -95 1015 -75
rect 15 -110 1015 -95
rect 15 -145 1015 -130
rect 15 -165 30 -145
rect 65 -165 85 -145
rect 105 -165 125 -145
rect 145 -165 165 -145
rect 185 -165 205 -145
rect 225 -165 245 -145
rect 265 -165 285 -145
rect 305 -165 325 -145
rect 345 -165 365 -145
rect 385 -165 405 -145
rect 425 -165 445 -145
rect 465 -165 485 -145
rect 505 -165 525 -145
rect 545 -165 565 -145
rect 585 -165 605 -145
rect 625 -165 645 -145
rect 665 -165 685 -145
rect 705 -165 725 -145
rect 745 -165 765 -145
rect 785 -165 805 -145
rect 825 -165 845 -145
rect 865 -165 885 -145
rect 905 -165 925 -145
rect 945 -165 965 -145
rect 1000 -165 1015 -145
rect 15 -180 1015 -165
rect 15 -215 1015 -200
rect 15 -235 30 -215
rect 65 -235 85 -215
rect 105 -235 125 -215
rect 145 -235 165 -215
rect 185 -235 205 -215
rect 225 -235 245 -215
rect 265 -235 285 -215
rect 305 -235 325 -215
rect 345 -235 365 -215
rect 385 -235 405 -215
rect 425 -235 445 -215
rect 465 -235 485 -215
rect 505 -235 525 -215
rect 545 -235 565 -215
rect 585 -235 605 -215
rect 625 -235 645 -215
rect 665 -235 685 -215
rect 705 -235 725 -215
rect 745 -235 765 -215
rect 785 -235 805 -215
rect 825 -235 845 -215
rect 865 -235 885 -215
rect 905 -235 925 -215
rect 945 -235 965 -215
rect 1000 -235 1015 -215
rect 15 -250 1015 -235
rect 15 -285 1015 -270
rect 15 -305 30 -285
rect 65 -305 85 -285
rect 105 -305 125 -285
rect 145 -305 165 -285
rect 185 -305 205 -285
rect 225 -305 245 -285
rect 265 -305 285 -285
rect 305 -305 325 -285
rect 345 -305 365 -285
rect 385 -305 405 -285
rect 425 -305 445 -285
rect 465 -305 485 -285
rect 505 -305 525 -285
rect 545 -305 565 -285
rect 585 -305 605 -285
rect 625 -305 645 -285
rect 665 -305 685 -285
rect 705 -305 725 -285
rect 745 -305 765 -285
rect 785 -305 805 -285
rect 825 -305 845 -285
rect 865 -305 885 -285
rect 905 -305 925 -285
rect 945 -305 965 -285
rect 1000 -305 1015 -285
rect 15 -320 1015 -305
rect 15 -355 1015 -340
rect 15 -375 30 -355
rect 65 -375 85 -355
rect 105 -375 125 -355
rect 145 -375 165 -355
rect 185 -375 205 -355
rect 225 -375 245 -355
rect 265 -375 285 -355
rect 305 -375 325 -355
rect 345 -375 365 -355
rect 385 -375 405 -355
rect 425 -375 445 -355
rect 465 -375 485 -355
rect 505 -375 525 -355
rect 545 -375 565 -355
rect 585 -375 605 -355
rect 625 -375 645 -355
rect 665 -375 685 -355
rect 705 -375 725 -355
rect 745 -375 765 -355
rect 785 -375 805 -355
rect 825 -375 845 -355
rect 865 -375 885 -355
rect 905 -375 925 -355
rect 945 -375 965 -355
rect 1000 -375 1015 -355
rect 15 -390 1015 -375
rect 15 -425 1015 -410
rect 15 -445 30 -425
rect 65 -445 85 -425
rect 105 -445 125 -425
rect 145 -445 165 -425
rect 185 -445 205 -425
rect 225 -445 245 -425
rect 265 -445 285 -425
rect 305 -445 325 -425
rect 345 -445 365 -425
rect 385 -445 405 -425
rect 425 -445 445 -425
rect 465 -445 485 -425
rect 505 -445 525 -425
rect 545 -445 565 -425
rect 585 -445 605 -425
rect 625 -445 645 -425
rect 665 -445 685 -425
rect 705 -445 725 -425
rect 745 -445 765 -425
rect 785 -445 805 -425
rect 825 -445 845 -425
rect 865 -445 885 -425
rect 905 -445 925 -425
rect 945 -445 965 -425
rect 1000 -445 1015 -425
rect 15 -460 1015 -445
rect 15 -495 1015 -480
rect 15 -515 30 -495
rect 65 -515 85 -495
rect 105 -515 125 -495
rect 145 -515 165 -495
rect 185 -515 205 -495
rect 225 -515 245 -495
rect 265 -515 285 -495
rect 305 -515 325 -495
rect 345 -515 365 -495
rect 385 -515 405 -495
rect 425 -515 445 -495
rect 465 -515 485 -495
rect 505 -515 525 -495
rect 545 -515 565 -495
rect 585 -515 605 -495
rect 625 -515 645 -495
rect 665 -515 685 -495
rect 705 -515 725 -495
rect 745 -515 765 -495
rect 785 -515 805 -495
rect 825 -515 845 -495
rect 865 -515 885 -495
rect 905 -515 925 -495
rect 945 -515 965 -495
rect 1000 -515 1015 -495
rect 15 -530 1015 -515
rect 15 -565 1015 -550
rect 15 -585 30 -565
rect 65 -585 85 -565
rect 105 -585 125 -565
rect 145 -585 165 -565
rect 185 -585 205 -565
rect 225 -585 245 -565
rect 265 -585 285 -565
rect 305 -585 325 -565
rect 345 -585 365 -565
rect 385 -585 405 -565
rect 425 -585 445 -565
rect 465 -585 485 -565
rect 505 -585 525 -565
rect 545 -585 565 -565
rect 585 -585 605 -565
rect 625 -585 645 -565
rect 665 -585 685 -565
rect 705 -585 725 -565
rect 745 -585 765 -565
rect 785 -585 805 -565
rect 825 -585 845 -565
rect 865 -585 885 -565
rect 905 -585 925 -565
rect 945 -585 965 -565
rect 1000 -585 1015 -565
rect 15 -595 1015 -585
rect -135 -675 1165 -665
rect -135 -695 -120 -675
rect -95 -695 -75 -675
rect -55 -695 -35 -675
rect -15 -695 5 -675
rect 25 -695 45 -675
rect 65 -695 85 -675
rect 105 -695 125 -675
rect 145 -695 165 -675
rect 185 -695 205 -675
rect 225 -695 245 -675
rect 265 -695 285 -675
rect 305 -695 325 -675
rect 345 -695 365 -675
rect 385 -695 405 -675
rect 425 -695 445 -675
rect 465 -695 485 -675
rect 505 -695 525 -675
rect 545 -695 565 -675
rect 585 -695 605 -675
rect 625 -695 645 -675
rect 665 -695 685 -675
rect 705 -695 725 -675
rect 745 -695 765 -675
rect 785 -695 805 -675
rect 825 -695 845 -675
rect 865 -695 885 -675
rect 905 -695 925 -675
rect 945 -695 965 -675
rect 985 -695 1005 -675
rect 1025 -695 1045 -675
rect 1065 -695 1085 -675
rect 1105 -695 1125 -675
rect 1150 -695 1165 -675
rect -135 -710 1165 -695
rect -135 -775 1165 -760
rect -135 -795 -120 -775
rect -95 -795 -75 -775
rect -55 -795 -35 -775
rect -15 -795 5 -775
rect 25 -795 45 -775
rect 65 -795 85 -775
rect 105 -795 125 -775
rect 145 -795 165 -775
rect 185 -795 205 -775
rect 225 -795 245 -775
rect 265 -795 285 -775
rect 305 -795 325 -775
rect 345 -795 365 -775
rect 385 -795 405 -775
rect 425 -795 445 -775
rect 465 -795 485 -775
rect 505 -795 525 -775
rect 545 -795 565 -775
rect 585 -795 605 -775
rect 625 -795 645 -775
rect 665 -795 685 -775
rect 705 -795 725 -775
rect 745 -795 765 -775
rect 785 -795 805 -775
rect 825 -795 845 -775
rect 865 -795 885 -775
rect 905 -795 925 -775
rect 945 -795 965 -775
rect 985 -795 1005 -775
rect 1025 -795 1045 -775
rect 1065 -795 1085 -775
rect 1105 -795 1125 -775
rect 1150 -795 1165 -775
rect -135 -810 1165 -795
rect -135 -875 1165 -860
rect -135 -895 -120 -875
rect -95 -895 -75 -875
rect -55 -895 -35 -875
rect -15 -895 5 -875
rect 25 -895 45 -875
rect 65 -895 85 -875
rect 105 -895 125 -875
rect 145 -895 165 -875
rect 185 -895 205 -875
rect 225 -895 245 -875
rect 265 -895 285 -875
rect 305 -895 325 -875
rect 345 -895 365 -875
rect 385 -895 405 -875
rect 425 -895 445 -875
rect 465 -895 485 -875
rect 505 -895 525 -875
rect 545 -895 565 -875
rect 585 -895 605 -875
rect 625 -895 645 -875
rect 665 -895 685 -875
rect 705 -895 725 -875
rect 745 -895 765 -875
rect 785 -895 805 -875
rect 825 -895 845 -875
rect 865 -895 885 -875
rect 905 -895 925 -875
rect 945 -895 965 -875
rect 985 -895 1005 -875
rect 1025 -895 1045 -875
rect 1065 -895 1085 -875
rect 1105 -895 1125 -875
rect 1150 -895 1165 -875
rect -135 -910 1165 -895
rect -135 -975 1165 -960
rect -135 -995 -120 -975
rect -95 -995 -75 -975
rect -55 -995 -35 -975
rect -15 -995 5 -975
rect 25 -995 45 -975
rect 65 -995 85 -975
rect 105 -995 125 -975
rect 145 -995 165 -975
rect 185 -995 205 -975
rect 225 -995 245 -975
rect 265 -995 285 -975
rect 305 -995 325 -975
rect 345 -995 365 -975
rect 385 -995 405 -975
rect 425 -995 445 -975
rect 465 -995 485 -975
rect 505 -995 525 -975
rect 545 -995 565 -975
rect 585 -995 605 -975
rect 625 -995 645 -975
rect 665 -995 685 -975
rect 705 -995 725 -975
rect 745 -995 765 -975
rect 785 -995 805 -975
rect 825 -995 845 -975
rect 865 -995 885 -975
rect 905 -995 925 -975
rect 945 -995 965 -975
rect 985 -995 1005 -975
rect 1025 -995 1045 -975
rect 1065 -995 1085 -975
rect 1105 -995 1125 -975
rect 1150 -995 1165 -975
rect -135 -1010 1165 -995
rect -135 -1075 1165 -1060
rect -135 -1095 -120 -1075
rect -95 -1095 -75 -1075
rect -55 -1095 -35 -1075
rect -15 -1095 5 -1075
rect 25 -1095 45 -1075
rect 65 -1095 85 -1075
rect 105 -1095 125 -1075
rect 145 -1095 165 -1075
rect 185 -1095 205 -1075
rect 225 -1095 245 -1075
rect 265 -1095 285 -1075
rect 305 -1095 325 -1075
rect 345 -1095 365 -1075
rect 385 -1095 405 -1075
rect 425 -1095 445 -1075
rect 465 -1095 485 -1075
rect 505 -1095 525 -1075
rect 545 -1095 565 -1075
rect 585 -1095 605 -1075
rect 625 -1095 645 -1075
rect 665 -1095 685 -1075
rect 705 -1095 725 -1075
rect 745 -1095 765 -1075
rect 785 -1095 805 -1075
rect 825 -1095 845 -1075
rect 865 -1095 885 -1075
rect 905 -1095 925 -1075
rect 945 -1095 965 -1075
rect 985 -1095 1005 -1075
rect 1025 -1095 1045 -1075
rect 1065 -1095 1085 -1075
rect 1105 -1095 1125 -1075
rect 1150 -1095 1165 -1075
rect -135 -1110 1165 -1095
rect -135 -1175 1165 -1160
rect -135 -1195 -120 -1175
rect -95 -1195 -75 -1175
rect -55 -1195 -35 -1175
rect -15 -1195 5 -1175
rect 25 -1195 45 -1175
rect 65 -1195 85 -1175
rect 105 -1195 125 -1175
rect 145 -1195 165 -1175
rect 185 -1195 205 -1175
rect 225 -1195 245 -1175
rect 265 -1195 285 -1175
rect 305 -1195 325 -1175
rect 345 -1195 365 -1175
rect 385 -1195 405 -1175
rect 425 -1195 445 -1175
rect 465 -1195 485 -1175
rect 505 -1195 525 -1175
rect 545 -1195 565 -1175
rect 585 -1195 605 -1175
rect 625 -1195 645 -1175
rect 665 -1195 685 -1175
rect 705 -1195 725 -1175
rect 745 -1195 765 -1175
rect 785 -1195 805 -1175
rect 825 -1195 845 -1175
rect 865 -1195 885 -1175
rect 905 -1195 925 -1175
rect 945 -1195 965 -1175
rect 985 -1195 1005 -1175
rect 1025 -1195 1045 -1175
rect 1065 -1195 1085 -1175
rect 1105 -1195 1125 -1175
rect 1150 -1195 1165 -1175
rect -135 -1205 1165 -1195
<< pdiff >>
rect -185 860 865 870
rect -185 840 -170 860
rect -135 840 -115 860
rect -95 840 -75 860
rect -55 840 -35 860
rect -15 840 5 860
rect 25 840 45 860
rect 65 840 85 860
rect 105 840 125 860
rect 145 840 165 860
rect 185 840 205 860
rect 225 840 245 860
rect 265 840 285 860
rect 305 840 325 860
rect 345 840 365 860
rect 385 840 405 860
rect 425 840 445 860
rect 465 840 485 860
rect 505 840 525 860
rect 545 840 565 860
rect 585 840 605 860
rect 625 840 645 860
rect 665 840 685 860
rect 705 840 725 860
rect 745 840 765 860
rect 785 840 805 860
rect 850 840 865 860
rect -185 825 865 840
rect -185 790 865 805
rect -185 770 -170 790
rect -135 770 -115 790
rect -95 770 -75 790
rect -55 770 -35 790
rect -15 770 5 790
rect 25 770 45 790
rect 65 770 85 790
rect 105 770 125 790
rect 145 770 165 790
rect 185 770 205 790
rect 225 770 245 790
rect 265 770 285 790
rect 305 770 325 790
rect 345 770 365 790
rect 385 770 405 790
rect 425 770 445 790
rect 465 770 485 790
rect 505 770 525 790
rect 545 770 565 790
rect 585 770 605 790
rect 625 770 645 790
rect 665 770 685 790
rect 705 770 725 790
rect 745 770 765 790
rect 785 770 805 790
rect 850 770 865 790
rect -185 755 865 770
rect -185 720 865 735
rect -185 700 -170 720
rect -135 700 -115 720
rect -95 700 -75 720
rect -55 700 -35 720
rect -15 700 5 720
rect 25 700 45 720
rect 65 700 85 720
rect 105 700 125 720
rect 145 700 165 720
rect 185 700 205 720
rect 225 700 245 720
rect 265 700 285 720
rect 305 700 325 720
rect 345 700 365 720
rect 385 700 405 720
rect 425 700 445 720
rect 465 700 485 720
rect 505 700 525 720
rect 545 700 565 720
rect 585 700 605 720
rect 625 700 645 720
rect 665 700 685 720
rect 705 700 725 720
rect 745 700 765 720
rect 785 700 805 720
rect 850 700 865 720
rect -185 685 865 700
rect -185 650 865 665
rect -185 630 -170 650
rect -135 630 -115 650
rect -95 630 -75 650
rect -55 630 -35 650
rect -15 630 5 650
rect 25 630 45 650
rect 65 630 85 650
rect 105 630 125 650
rect 145 630 165 650
rect 185 630 205 650
rect 225 630 245 650
rect 265 630 285 650
rect 305 630 325 650
rect 345 630 365 650
rect 385 630 405 650
rect 425 630 445 650
rect 465 630 485 650
rect 505 630 525 650
rect 545 630 565 650
rect 585 630 605 650
rect 625 630 645 650
rect 665 630 685 650
rect 705 630 725 650
rect 745 630 765 650
rect 785 630 805 650
rect 850 630 865 650
rect -185 615 865 630
rect -185 580 865 595
rect -185 560 -170 580
rect -135 560 -115 580
rect -95 560 -75 580
rect -55 560 -35 580
rect -15 560 5 580
rect 25 560 45 580
rect 65 560 85 580
rect 105 560 125 580
rect 145 560 165 580
rect 185 560 205 580
rect 225 560 245 580
rect 265 560 285 580
rect 305 560 325 580
rect 345 560 365 580
rect 385 560 405 580
rect 425 560 445 580
rect 465 560 485 580
rect 505 560 525 580
rect 545 560 565 580
rect 585 560 605 580
rect 625 560 645 580
rect 665 560 685 580
rect 705 560 725 580
rect 745 560 765 580
rect 785 560 805 580
rect 850 560 865 580
rect -185 550 865 560
<< ndiffc >>
rect 30 465 65 485
rect 85 465 105 485
rect 125 465 145 485
rect 165 465 185 485
rect 205 465 225 485
rect 245 465 265 485
rect 285 465 305 485
rect 325 465 345 485
rect 365 465 385 485
rect 405 465 425 485
rect 445 465 465 485
rect 485 465 505 485
rect 525 465 545 485
rect 565 465 585 485
rect 605 465 625 485
rect 645 465 665 485
rect 685 465 705 485
rect 725 465 745 485
rect 765 465 785 485
rect 805 465 825 485
rect 845 465 865 485
rect 885 465 905 485
rect 925 465 945 485
rect 965 465 1000 485
rect 30 395 65 415
rect 85 395 105 415
rect 125 395 145 415
rect 165 395 185 415
rect 205 395 225 415
rect 245 395 265 415
rect 285 395 305 415
rect 325 395 345 415
rect 365 395 385 415
rect 405 395 425 415
rect 445 395 465 415
rect 485 395 505 415
rect 525 395 545 415
rect 565 395 585 415
rect 605 395 625 415
rect 645 395 665 415
rect 685 395 705 415
rect 725 395 745 415
rect 765 395 785 415
rect 805 395 825 415
rect 845 395 865 415
rect 885 395 905 415
rect 925 395 945 415
rect 965 395 1000 415
rect 30 325 65 345
rect 85 325 105 345
rect 125 325 145 345
rect 165 325 185 345
rect 205 325 225 345
rect 245 325 265 345
rect 285 325 305 345
rect 325 325 345 345
rect 365 325 385 345
rect 405 325 425 345
rect 445 325 465 345
rect 485 325 505 345
rect 525 325 545 345
rect 565 325 585 345
rect 605 325 625 345
rect 645 325 665 345
rect 685 325 705 345
rect 725 325 745 345
rect 765 325 785 345
rect 805 325 825 345
rect 845 325 865 345
rect 885 325 905 345
rect 925 325 945 345
rect 965 325 1000 345
rect 30 255 65 275
rect 85 255 105 275
rect 125 255 145 275
rect 165 255 185 275
rect 205 255 225 275
rect 245 255 265 275
rect 285 255 305 275
rect 325 255 345 275
rect 365 255 385 275
rect 405 255 425 275
rect 445 255 465 275
rect 485 255 505 275
rect 525 255 545 275
rect 565 255 585 275
rect 605 255 625 275
rect 645 255 665 275
rect 685 255 705 275
rect 725 255 745 275
rect 765 255 785 275
rect 805 255 825 275
rect 845 255 865 275
rect 885 255 905 275
rect 925 255 945 275
rect 965 255 1000 275
rect 30 185 65 205
rect 85 185 105 205
rect 125 185 145 205
rect 165 185 185 205
rect 205 185 225 205
rect 245 185 265 205
rect 285 185 305 205
rect 325 185 345 205
rect 365 185 385 205
rect 405 185 425 205
rect 445 185 465 205
rect 485 185 505 205
rect 525 185 545 205
rect 565 185 585 205
rect 605 185 625 205
rect 645 185 665 205
rect 685 185 705 205
rect 725 185 745 205
rect 765 185 785 205
rect 805 185 825 205
rect 845 185 865 205
rect 885 185 905 205
rect 925 185 945 205
rect 965 185 1000 205
rect 30 115 65 135
rect 85 115 105 135
rect 125 115 145 135
rect 165 115 185 135
rect 205 115 225 135
rect 245 115 265 135
rect 285 115 305 135
rect 325 115 345 135
rect 365 115 385 135
rect 405 115 425 135
rect 445 115 465 135
rect 485 115 505 135
rect 525 115 545 135
rect 565 115 585 135
rect 605 115 625 135
rect 645 115 665 135
rect 685 115 705 135
rect 725 115 745 135
rect 765 115 785 135
rect 805 115 825 135
rect 845 115 865 135
rect 885 115 905 135
rect 925 115 945 135
rect 965 115 1000 135
rect 30 45 65 65
rect 85 45 105 65
rect 125 45 145 65
rect 165 45 185 65
rect 205 45 225 65
rect 245 45 265 65
rect 285 45 305 65
rect 325 45 345 65
rect 365 45 385 65
rect 405 45 425 65
rect 445 45 465 65
rect 485 45 505 65
rect 525 45 545 65
rect 565 45 585 65
rect 605 45 625 65
rect 645 45 665 65
rect 685 45 705 65
rect 725 45 745 65
rect 765 45 785 65
rect 805 45 825 65
rect 845 45 865 65
rect 885 45 905 65
rect 925 45 945 65
rect 965 45 1000 65
rect 30 -25 65 -5
rect 85 -25 105 -5
rect 125 -25 145 -5
rect 165 -25 185 -5
rect 205 -25 225 -5
rect 245 -25 265 -5
rect 285 -25 305 -5
rect 325 -25 345 -5
rect 365 -25 385 -5
rect 405 -25 425 -5
rect 445 -25 465 -5
rect 485 -25 505 -5
rect 525 -25 545 -5
rect 565 -25 585 -5
rect 605 -25 625 -5
rect 645 -25 665 -5
rect 685 -25 705 -5
rect 725 -25 745 -5
rect 765 -25 785 -5
rect 805 -25 825 -5
rect 845 -25 865 -5
rect 885 -25 905 -5
rect 925 -25 945 -5
rect 965 -25 1000 -5
rect 30 -95 65 -75
rect 85 -95 105 -75
rect 125 -95 145 -75
rect 165 -95 185 -75
rect 205 -95 225 -75
rect 245 -95 265 -75
rect 285 -95 305 -75
rect 325 -95 345 -75
rect 365 -95 385 -75
rect 405 -95 425 -75
rect 445 -95 465 -75
rect 485 -95 505 -75
rect 525 -95 545 -75
rect 565 -95 585 -75
rect 605 -95 625 -75
rect 645 -95 665 -75
rect 685 -95 705 -75
rect 725 -95 745 -75
rect 765 -95 785 -75
rect 805 -95 825 -75
rect 845 -95 865 -75
rect 885 -95 905 -75
rect 925 -95 945 -75
rect 965 -95 1000 -75
rect 30 -165 65 -145
rect 85 -165 105 -145
rect 125 -165 145 -145
rect 165 -165 185 -145
rect 205 -165 225 -145
rect 245 -165 265 -145
rect 285 -165 305 -145
rect 325 -165 345 -145
rect 365 -165 385 -145
rect 405 -165 425 -145
rect 445 -165 465 -145
rect 485 -165 505 -145
rect 525 -165 545 -145
rect 565 -165 585 -145
rect 605 -165 625 -145
rect 645 -165 665 -145
rect 685 -165 705 -145
rect 725 -165 745 -145
rect 765 -165 785 -145
rect 805 -165 825 -145
rect 845 -165 865 -145
rect 885 -165 905 -145
rect 925 -165 945 -145
rect 965 -165 1000 -145
rect 30 -235 65 -215
rect 85 -235 105 -215
rect 125 -235 145 -215
rect 165 -235 185 -215
rect 205 -235 225 -215
rect 245 -235 265 -215
rect 285 -235 305 -215
rect 325 -235 345 -215
rect 365 -235 385 -215
rect 405 -235 425 -215
rect 445 -235 465 -215
rect 485 -235 505 -215
rect 525 -235 545 -215
rect 565 -235 585 -215
rect 605 -235 625 -215
rect 645 -235 665 -215
rect 685 -235 705 -215
rect 725 -235 745 -215
rect 765 -235 785 -215
rect 805 -235 825 -215
rect 845 -235 865 -215
rect 885 -235 905 -215
rect 925 -235 945 -215
rect 965 -235 1000 -215
rect 30 -305 65 -285
rect 85 -305 105 -285
rect 125 -305 145 -285
rect 165 -305 185 -285
rect 205 -305 225 -285
rect 245 -305 265 -285
rect 285 -305 305 -285
rect 325 -305 345 -285
rect 365 -305 385 -285
rect 405 -305 425 -285
rect 445 -305 465 -285
rect 485 -305 505 -285
rect 525 -305 545 -285
rect 565 -305 585 -285
rect 605 -305 625 -285
rect 645 -305 665 -285
rect 685 -305 705 -285
rect 725 -305 745 -285
rect 765 -305 785 -285
rect 805 -305 825 -285
rect 845 -305 865 -285
rect 885 -305 905 -285
rect 925 -305 945 -285
rect 965 -305 1000 -285
rect 30 -375 65 -355
rect 85 -375 105 -355
rect 125 -375 145 -355
rect 165 -375 185 -355
rect 205 -375 225 -355
rect 245 -375 265 -355
rect 285 -375 305 -355
rect 325 -375 345 -355
rect 365 -375 385 -355
rect 405 -375 425 -355
rect 445 -375 465 -355
rect 485 -375 505 -355
rect 525 -375 545 -355
rect 565 -375 585 -355
rect 605 -375 625 -355
rect 645 -375 665 -355
rect 685 -375 705 -355
rect 725 -375 745 -355
rect 765 -375 785 -355
rect 805 -375 825 -355
rect 845 -375 865 -355
rect 885 -375 905 -355
rect 925 -375 945 -355
rect 965 -375 1000 -355
rect 30 -445 65 -425
rect 85 -445 105 -425
rect 125 -445 145 -425
rect 165 -445 185 -425
rect 205 -445 225 -425
rect 245 -445 265 -425
rect 285 -445 305 -425
rect 325 -445 345 -425
rect 365 -445 385 -425
rect 405 -445 425 -425
rect 445 -445 465 -425
rect 485 -445 505 -425
rect 525 -445 545 -425
rect 565 -445 585 -425
rect 605 -445 625 -425
rect 645 -445 665 -425
rect 685 -445 705 -425
rect 725 -445 745 -425
rect 765 -445 785 -425
rect 805 -445 825 -425
rect 845 -445 865 -425
rect 885 -445 905 -425
rect 925 -445 945 -425
rect 965 -445 1000 -425
rect 30 -515 65 -495
rect 85 -515 105 -495
rect 125 -515 145 -495
rect 165 -515 185 -495
rect 205 -515 225 -495
rect 245 -515 265 -495
rect 285 -515 305 -495
rect 325 -515 345 -495
rect 365 -515 385 -495
rect 405 -515 425 -495
rect 445 -515 465 -495
rect 485 -515 505 -495
rect 525 -515 545 -495
rect 565 -515 585 -495
rect 605 -515 625 -495
rect 645 -515 665 -495
rect 685 -515 705 -495
rect 725 -515 745 -495
rect 765 -515 785 -495
rect 805 -515 825 -495
rect 845 -515 865 -495
rect 885 -515 905 -495
rect 925 -515 945 -495
rect 965 -515 1000 -495
rect 30 -585 65 -565
rect 85 -585 105 -565
rect 125 -585 145 -565
rect 165 -585 185 -565
rect 205 -585 225 -565
rect 245 -585 265 -565
rect 285 -585 305 -565
rect 325 -585 345 -565
rect 365 -585 385 -565
rect 405 -585 425 -565
rect 445 -585 465 -565
rect 485 -585 505 -565
rect 525 -585 545 -565
rect 565 -585 585 -565
rect 605 -585 625 -565
rect 645 -585 665 -565
rect 685 -585 705 -565
rect 725 -585 745 -565
rect 765 -585 785 -565
rect 805 -585 825 -565
rect 845 -585 865 -565
rect 885 -585 905 -565
rect 925 -585 945 -565
rect 965 -585 1000 -565
rect -120 -695 -95 -675
rect -75 -695 -55 -675
rect -35 -695 -15 -675
rect 5 -695 25 -675
rect 45 -695 65 -675
rect 85 -695 105 -675
rect 125 -695 145 -675
rect 165 -695 185 -675
rect 205 -695 225 -675
rect 245 -695 265 -675
rect 285 -695 305 -675
rect 325 -695 345 -675
rect 365 -695 385 -675
rect 405 -695 425 -675
rect 445 -695 465 -675
rect 485 -695 505 -675
rect 525 -695 545 -675
rect 565 -695 585 -675
rect 605 -695 625 -675
rect 645 -695 665 -675
rect 685 -695 705 -675
rect 725 -695 745 -675
rect 765 -695 785 -675
rect 805 -695 825 -675
rect 845 -695 865 -675
rect 885 -695 905 -675
rect 925 -695 945 -675
rect 965 -695 985 -675
rect 1005 -695 1025 -675
rect 1045 -695 1065 -675
rect 1085 -695 1105 -675
rect 1125 -695 1150 -675
rect -120 -795 -95 -775
rect -75 -795 -55 -775
rect -35 -795 -15 -775
rect 5 -795 25 -775
rect 45 -795 65 -775
rect 85 -795 105 -775
rect 125 -795 145 -775
rect 165 -795 185 -775
rect 205 -795 225 -775
rect 245 -795 265 -775
rect 285 -795 305 -775
rect 325 -795 345 -775
rect 365 -795 385 -775
rect 405 -795 425 -775
rect 445 -795 465 -775
rect 485 -795 505 -775
rect 525 -795 545 -775
rect 565 -795 585 -775
rect 605 -795 625 -775
rect 645 -795 665 -775
rect 685 -795 705 -775
rect 725 -795 745 -775
rect 765 -795 785 -775
rect 805 -795 825 -775
rect 845 -795 865 -775
rect 885 -795 905 -775
rect 925 -795 945 -775
rect 965 -795 985 -775
rect 1005 -795 1025 -775
rect 1045 -795 1065 -775
rect 1085 -795 1105 -775
rect 1125 -795 1150 -775
rect -120 -895 -95 -875
rect -75 -895 -55 -875
rect -35 -895 -15 -875
rect 5 -895 25 -875
rect 45 -895 65 -875
rect 85 -895 105 -875
rect 125 -895 145 -875
rect 165 -895 185 -875
rect 205 -895 225 -875
rect 245 -895 265 -875
rect 285 -895 305 -875
rect 325 -895 345 -875
rect 365 -895 385 -875
rect 405 -895 425 -875
rect 445 -895 465 -875
rect 485 -895 505 -875
rect 525 -895 545 -875
rect 565 -895 585 -875
rect 605 -895 625 -875
rect 645 -895 665 -875
rect 685 -895 705 -875
rect 725 -895 745 -875
rect 765 -895 785 -875
rect 805 -895 825 -875
rect 845 -895 865 -875
rect 885 -895 905 -875
rect 925 -895 945 -875
rect 965 -895 985 -875
rect 1005 -895 1025 -875
rect 1045 -895 1065 -875
rect 1085 -895 1105 -875
rect 1125 -895 1150 -875
rect -120 -995 -95 -975
rect -75 -995 -55 -975
rect -35 -995 -15 -975
rect 5 -995 25 -975
rect 45 -995 65 -975
rect 85 -995 105 -975
rect 125 -995 145 -975
rect 165 -995 185 -975
rect 205 -995 225 -975
rect 245 -995 265 -975
rect 285 -995 305 -975
rect 325 -995 345 -975
rect 365 -995 385 -975
rect 405 -995 425 -975
rect 445 -995 465 -975
rect 485 -995 505 -975
rect 525 -995 545 -975
rect 565 -995 585 -975
rect 605 -995 625 -975
rect 645 -995 665 -975
rect 685 -995 705 -975
rect 725 -995 745 -975
rect 765 -995 785 -975
rect 805 -995 825 -975
rect 845 -995 865 -975
rect 885 -995 905 -975
rect 925 -995 945 -975
rect 965 -995 985 -975
rect 1005 -995 1025 -975
rect 1045 -995 1065 -975
rect 1085 -995 1105 -975
rect 1125 -995 1150 -975
rect -120 -1095 -95 -1075
rect -75 -1095 -55 -1075
rect -35 -1095 -15 -1075
rect 5 -1095 25 -1075
rect 45 -1095 65 -1075
rect 85 -1095 105 -1075
rect 125 -1095 145 -1075
rect 165 -1095 185 -1075
rect 205 -1095 225 -1075
rect 245 -1095 265 -1075
rect 285 -1095 305 -1075
rect 325 -1095 345 -1075
rect 365 -1095 385 -1075
rect 405 -1095 425 -1075
rect 445 -1095 465 -1075
rect 485 -1095 505 -1075
rect 525 -1095 545 -1075
rect 565 -1095 585 -1075
rect 605 -1095 625 -1075
rect 645 -1095 665 -1075
rect 685 -1095 705 -1075
rect 725 -1095 745 -1075
rect 765 -1095 785 -1075
rect 805 -1095 825 -1075
rect 845 -1095 865 -1075
rect 885 -1095 905 -1075
rect 925 -1095 945 -1075
rect 965 -1095 985 -1075
rect 1005 -1095 1025 -1075
rect 1045 -1095 1065 -1075
rect 1085 -1095 1105 -1075
rect 1125 -1095 1150 -1075
rect -120 -1195 -95 -1175
rect -75 -1195 -55 -1175
rect -35 -1195 -15 -1175
rect 5 -1195 25 -1175
rect 45 -1195 65 -1175
rect 85 -1195 105 -1175
rect 125 -1195 145 -1175
rect 165 -1195 185 -1175
rect 205 -1195 225 -1175
rect 245 -1195 265 -1175
rect 285 -1195 305 -1175
rect 325 -1195 345 -1175
rect 365 -1195 385 -1175
rect 405 -1195 425 -1175
rect 445 -1195 465 -1175
rect 485 -1195 505 -1175
rect 525 -1195 545 -1175
rect 565 -1195 585 -1175
rect 605 -1195 625 -1175
rect 645 -1195 665 -1175
rect 685 -1195 705 -1175
rect 725 -1195 745 -1175
rect 765 -1195 785 -1175
rect 805 -1195 825 -1175
rect 845 -1195 865 -1175
rect 885 -1195 905 -1175
rect 925 -1195 945 -1175
rect 965 -1195 985 -1175
rect 1005 -1195 1025 -1175
rect 1045 -1195 1065 -1175
rect 1085 -1195 1105 -1175
rect 1125 -1195 1150 -1175
<< pdiffc >>
rect -170 840 -135 860
rect -115 840 -95 860
rect -75 840 -55 860
rect -35 840 -15 860
rect 5 840 25 860
rect 45 840 65 860
rect 85 840 105 860
rect 125 840 145 860
rect 165 840 185 860
rect 205 840 225 860
rect 245 840 265 860
rect 285 840 305 860
rect 325 840 345 860
rect 365 840 385 860
rect 405 840 425 860
rect 445 840 465 860
rect 485 840 505 860
rect 525 840 545 860
rect 565 840 585 860
rect 605 840 625 860
rect 645 840 665 860
rect 685 840 705 860
rect 725 840 745 860
rect 765 840 785 860
rect 805 840 850 860
rect -170 770 -135 790
rect -115 770 -95 790
rect -75 770 -55 790
rect -35 770 -15 790
rect 5 770 25 790
rect 45 770 65 790
rect 85 770 105 790
rect 125 770 145 790
rect 165 770 185 790
rect 205 770 225 790
rect 245 770 265 790
rect 285 770 305 790
rect 325 770 345 790
rect 365 770 385 790
rect 405 770 425 790
rect 445 770 465 790
rect 485 770 505 790
rect 525 770 545 790
rect 565 770 585 790
rect 605 770 625 790
rect 645 770 665 790
rect 685 770 705 790
rect 725 770 745 790
rect 765 770 785 790
rect 805 770 850 790
rect -170 700 -135 720
rect -115 700 -95 720
rect -75 700 -55 720
rect -35 700 -15 720
rect 5 700 25 720
rect 45 700 65 720
rect 85 700 105 720
rect 125 700 145 720
rect 165 700 185 720
rect 205 700 225 720
rect 245 700 265 720
rect 285 700 305 720
rect 325 700 345 720
rect 365 700 385 720
rect 405 700 425 720
rect 445 700 465 720
rect 485 700 505 720
rect 525 700 545 720
rect 565 700 585 720
rect 605 700 625 720
rect 645 700 665 720
rect 685 700 705 720
rect 725 700 745 720
rect 765 700 785 720
rect 805 700 850 720
rect -170 630 -135 650
rect -115 630 -95 650
rect -75 630 -55 650
rect -35 630 -15 650
rect 5 630 25 650
rect 45 630 65 650
rect 85 630 105 650
rect 125 630 145 650
rect 165 630 185 650
rect 205 630 225 650
rect 245 630 265 650
rect 285 630 305 650
rect 325 630 345 650
rect 365 630 385 650
rect 405 630 425 650
rect 445 630 465 650
rect 485 630 505 650
rect 525 630 545 650
rect 565 630 585 650
rect 605 630 625 650
rect 645 630 665 650
rect 685 630 705 650
rect 725 630 745 650
rect 765 630 785 650
rect 805 630 850 650
rect -170 560 -135 580
rect -115 560 -95 580
rect -75 560 -55 580
rect -35 560 -15 580
rect 5 560 25 580
rect 45 560 65 580
rect 85 560 105 580
rect 125 560 145 580
rect 165 560 185 580
rect 205 560 225 580
rect 245 560 265 580
rect 285 560 305 580
rect 325 560 345 580
rect 365 560 385 580
rect 405 560 425 580
rect 445 560 465 580
rect 485 560 505 580
rect 525 560 545 580
rect 565 560 585 580
rect 605 560 625 580
rect 645 560 665 580
rect 685 560 705 580
rect 725 560 745 580
rect 765 560 785 580
rect 805 560 850 580
<< psubdiff >>
rect -135 -635 1165 -625
rect -135 -655 -120 -635
rect -95 -655 -75 -635
rect -55 -655 -35 -635
rect -15 -655 5 -635
rect 25 -655 45 -635
rect 65 -655 85 -635
rect 105 -655 125 -635
rect 145 -655 165 -635
rect 185 -655 205 -635
rect 225 -655 245 -635
rect 265 -655 285 -635
rect 305 -655 325 -635
rect 345 -655 365 -635
rect 385 -655 405 -635
rect 425 -655 445 -635
rect 465 -655 485 -635
rect 505 -655 525 -635
rect 545 -655 565 -635
rect 585 -655 605 -635
rect 625 -655 645 -635
rect 665 -655 685 -635
rect 705 -655 725 -635
rect 745 -655 765 -635
rect 785 -655 805 -635
rect 825 -655 845 -635
rect 865 -655 885 -635
rect 905 -655 925 -635
rect 945 -655 965 -635
rect 985 -655 1005 -635
rect 1025 -655 1045 -635
rect 1065 -655 1085 -635
rect 1105 -655 1125 -635
rect 1150 -655 1165 -635
rect -135 -665 1165 -655
<< nsubdiff >>
rect -185 900 865 910
rect -185 880 -170 900
rect -135 880 -115 900
rect -95 880 -75 900
rect -55 880 -35 900
rect -15 880 5 900
rect 25 880 45 900
rect 65 880 85 900
rect 105 880 125 900
rect 145 880 165 900
rect 185 880 205 900
rect 225 880 245 900
rect 265 880 285 900
rect 305 880 325 900
rect 345 880 365 900
rect 385 880 405 900
rect 425 880 445 900
rect 465 880 485 900
rect 505 880 525 900
rect 545 880 565 900
rect 585 880 605 900
rect 625 880 645 900
rect 665 880 685 900
rect 705 880 725 900
rect 745 880 765 900
rect 785 880 805 900
rect 850 880 865 900
rect -185 870 865 880
<< psubdiffcont >>
rect -120 -655 -95 -635
rect -75 -655 -55 -635
rect -35 -655 -15 -635
rect 5 -655 25 -635
rect 45 -655 65 -635
rect 85 -655 105 -635
rect 125 -655 145 -635
rect 165 -655 185 -635
rect 205 -655 225 -635
rect 245 -655 265 -635
rect 285 -655 305 -635
rect 325 -655 345 -635
rect 365 -655 385 -635
rect 405 -655 425 -635
rect 445 -655 465 -635
rect 485 -655 505 -635
rect 525 -655 545 -635
rect 565 -655 585 -635
rect 605 -655 625 -635
rect 645 -655 665 -635
rect 685 -655 705 -635
rect 725 -655 745 -635
rect 765 -655 785 -635
rect 805 -655 825 -635
rect 845 -655 865 -635
rect 885 -655 905 -635
rect 925 -655 945 -635
rect 965 -655 985 -635
rect 1005 -655 1025 -635
rect 1045 -655 1065 -635
rect 1085 -655 1105 -635
rect 1125 -655 1150 -635
<< nsubdiffcont >>
rect -170 880 -135 900
rect -115 880 -95 900
rect -75 880 -55 900
rect -35 880 -15 900
rect 5 880 25 900
rect 45 880 65 900
rect 85 880 105 900
rect 125 880 145 900
rect 165 880 185 900
rect 205 880 225 900
rect 245 880 265 900
rect 285 880 305 900
rect 325 880 345 900
rect 365 880 385 900
rect 405 880 425 900
rect 445 880 465 900
rect 485 880 505 900
rect 525 880 545 900
rect 565 880 585 900
rect 605 880 625 900
rect 645 880 665 900
rect 685 880 705 900
rect 725 880 745 900
rect 765 880 785 900
rect 805 880 850 900
<< poly >>
rect -215 805 -185 825
rect 865 805 880 825
rect -215 755 -200 805
rect -215 735 -185 755
rect 865 735 880 755
rect -215 685 -200 735
rect -215 665 -185 685
rect 865 665 880 685
rect -215 615 -200 665
rect -215 595 -185 615
rect 865 595 880 615
rect 1025 450 1190 460
rect 0 430 15 450
rect 1015 430 1035 450
rect 1060 430 1080 450
rect 1100 430 1120 450
rect 1140 430 1160 450
rect 1180 430 1190 450
rect 1025 420 1190 430
rect 1025 380 1190 390
rect 0 360 15 380
rect 1015 360 1035 380
rect 1060 360 1080 380
rect 1100 360 1120 380
rect 1140 360 1160 380
rect 1180 360 1190 380
rect 1025 350 1190 360
rect 1025 310 1190 320
rect 0 290 15 310
rect 1015 290 1035 310
rect 1060 290 1080 310
rect 1100 290 1120 310
rect 1140 290 1160 310
rect 1180 290 1190 310
rect 1025 280 1190 290
rect 1025 240 1190 250
rect 0 220 15 240
rect 1015 220 1035 240
rect 1060 220 1080 240
rect 1100 220 1120 240
rect 1140 220 1160 240
rect 1180 220 1190 240
rect 1025 210 1190 220
rect 1025 170 1190 180
rect 0 150 15 170
rect 1015 150 1035 170
rect 1060 150 1080 170
rect 1100 150 1120 170
rect 1140 150 1160 170
rect 1180 150 1190 170
rect 1025 140 1190 150
rect 1025 100 1190 110
rect 0 80 15 100
rect 1015 80 1035 100
rect 1060 80 1080 100
rect 1100 80 1120 100
rect 1140 80 1160 100
rect 1180 80 1190 100
rect 1025 70 1190 80
rect 1025 30 1190 40
rect 0 10 15 30
rect 1015 10 1035 30
rect 1060 10 1080 30
rect 1100 10 1120 30
rect 1140 10 1160 30
rect 1180 10 1190 30
rect 1025 0 1190 10
rect 1025 -40 1190 -30
rect 0 -60 15 -40
rect 1015 -60 1035 -40
rect 1060 -60 1080 -40
rect 1100 -60 1120 -40
rect 1140 -60 1160 -40
rect 1180 -60 1190 -40
rect 1025 -70 1190 -60
rect 1025 -110 1190 -100
rect 0 -130 15 -110
rect 1015 -130 1035 -110
rect 1060 -130 1080 -110
rect 1100 -130 1120 -110
rect 1140 -130 1160 -110
rect 1180 -130 1190 -110
rect 1025 -140 1190 -130
rect 1025 -180 1190 -170
rect 0 -200 15 -180
rect 1015 -200 1035 -180
rect 1060 -200 1080 -180
rect 1100 -200 1120 -180
rect 1140 -200 1160 -180
rect 1180 -200 1190 -180
rect 1025 -210 1190 -200
rect 1025 -250 1190 -240
rect 0 -270 15 -250
rect 1015 -270 1035 -250
rect 1060 -270 1080 -250
rect 1100 -270 1120 -250
rect 1140 -270 1160 -250
rect 1180 -270 1190 -250
rect 1025 -280 1190 -270
rect 1025 -320 1190 -310
rect 0 -340 15 -320
rect 1015 -340 1035 -320
rect 1060 -340 1080 -320
rect 1100 -340 1120 -320
rect 1140 -340 1160 -320
rect 1180 -340 1190 -320
rect 1025 -350 1190 -340
rect 1025 -390 1190 -380
rect 0 -410 15 -390
rect 1015 -410 1035 -390
rect 1060 -410 1080 -390
rect 1100 -410 1120 -390
rect 1140 -410 1160 -390
rect 1180 -410 1190 -390
rect 1025 -420 1190 -410
rect 1025 -460 1190 -450
rect 0 -480 15 -460
rect 1015 -480 1035 -460
rect 1060 -480 1080 -460
rect 1100 -480 1120 -460
rect 1140 -480 1160 -460
rect 1180 -480 1190 -460
rect 1025 -490 1190 -480
rect 1025 -530 1190 -520
rect 0 -550 15 -530
rect 1015 -550 1035 -530
rect 1060 -550 1080 -530
rect 1100 -550 1120 -530
rect 1140 -550 1160 -530
rect 1180 -550 1190 -530
rect 1025 -560 1190 -550
rect -310 -720 -135 -710
rect -310 -750 -300 -720
rect -280 -750 -260 -720
rect -240 -750 -220 -720
rect -200 -750 -180 -720
rect -155 -750 -135 -720
rect -310 -760 -135 -750
rect 1165 -760 1180 -710
rect -310 -820 -135 -810
rect -310 -850 -300 -820
rect -280 -850 -260 -820
rect -240 -850 -220 -820
rect -200 -850 -180 -820
rect -155 -850 -135 -820
rect -310 -860 -135 -850
rect 1165 -860 1180 -810
rect -310 -920 -135 -910
rect -310 -950 -300 -920
rect -280 -950 -260 -920
rect -240 -950 -220 -920
rect -200 -950 -180 -920
rect -155 -950 -135 -920
rect -310 -960 -135 -950
rect 1165 -960 1180 -910
rect -310 -1020 -135 -1010
rect -310 -1050 -300 -1020
rect -280 -1050 -260 -1020
rect -240 -1050 -220 -1020
rect -200 -1050 -180 -1020
rect -155 -1050 -135 -1020
rect -310 -1060 -135 -1050
rect 1165 -1060 1180 -1010
rect -310 -1120 -135 -1110
rect -310 -1150 -300 -1120
rect -280 -1150 -260 -1120
rect -240 -1150 -220 -1120
rect -200 -1150 -180 -1120
rect -155 -1150 -135 -1120
rect -310 -1160 -135 -1150
rect 1165 -1160 1180 -1110
<< polycont >>
rect 1035 430 1060 450
rect 1080 430 1100 450
rect 1120 430 1140 450
rect 1160 430 1180 450
rect 1035 360 1060 380
rect 1080 360 1100 380
rect 1120 360 1140 380
rect 1160 360 1180 380
rect 1035 290 1060 310
rect 1080 290 1100 310
rect 1120 290 1140 310
rect 1160 290 1180 310
rect 1035 220 1060 240
rect 1080 220 1100 240
rect 1120 220 1140 240
rect 1160 220 1180 240
rect 1035 150 1060 170
rect 1080 150 1100 170
rect 1120 150 1140 170
rect 1160 150 1180 170
rect 1035 80 1060 100
rect 1080 80 1100 100
rect 1120 80 1140 100
rect 1160 80 1180 100
rect 1035 10 1060 30
rect 1080 10 1100 30
rect 1120 10 1140 30
rect 1160 10 1180 30
rect 1035 -60 1060 -40
rect 1080 -60 1100 -40
rect 1120 -60 1140 -40
rect 1160 -60 1180 -40
rect 1035 -130 1060 -110
rect 1080 -130 1100 -110
rect 1120 -130 1140 -110
rect 1160 -130 1180 -110
rect 1035 -200 1060 -180
rect 1080 -200 1100 -180
rect 1120 -200 1140 -180
rect 1160 -200 1180 -180
rect 1035 -270 1060 -250
rect 1080 -270 1100 -250
rect 1120 -270 1140 -250
rect 1160 -270 1180 -250
rect 1035 -340 1060 -320
rect 1080 -340 1100 -320
rect 1120 -340 1140 -320
rect 1160 -340 1180 -320
rect 1035 -410 1060 -390
rect 1080 -410 1100 -390
rect 1120 -410 1140 -390
rect 1160 -410 1180 -390
rect 1035 -480 1060 -460
rect 1080 -480 1100 -460
rect 1120 -480 1140 -460
rect 1160 -480 1180 -460
rect 1035 -550 1060 -530
rect 1080 -550 1100 -530
rect 1120 -550 1140 -530
rect 1160 -550 1180 -530
rect -300 -750 -280 -720
rect -260 -750 -240 -720
rect -220 -750 -200 -720
rect -180 -750 -155 -720
rect -300 -850 -280 -820
rect -260 -850 -240 -820
rect -220 -850 -200 -820
rect -180 -850 -155 -820
rect -300 -950 -280 -920
rect -260 -950 -240 -920
rect -220 -950 -200 -920
rect -180 -950 -155 -920
rect -300 -1050 -280 -1020
rect -260 -1050 -240 -1020
rect -220 -1050 -200 -1020
rect -180 -1050 -155 -1020
rect -300 -1150 -280 -1120
rect -260 -1150 -240 -1120
rect -220 -1150 -200 -1120
rect -180 -1150 -155 -1120
<< locali >>
rect -185 900 865 910
rect -185 880 -170 900
rect -135 880 -115 900
rect -95 880 -75 900
rect -55 880 -35 900
rect -15 880 5 900
rect 25 880 45 900
rect 65 880 85 900
rect 105 880 125 900
rect 145 880 165 900
rect 185 880 205 900
rect 225 880 245 900
rect 265 880 285 900
rect 305 880 325 900
rect 345 880 365 900
rect 385 880 405 900
rect 425 880 445 900
rect 465 880 485 900
rect 505 880 525 900
rect 545 880 565 900
rect 585 880 605 900
rect 625 880 645 900
rect 665 880 685 900
rect 705 880 725 900
rect 745 880 765 900
rect 785 880 805 900
rect 850 880 865 900
rect -185 860 865 880
rect -185 840 -170 860
rect -135 840 -115 860
rect -95 840 -75 860
rect -55 840 -35 860
rect -15 840 5 860
rect 25 840 45 860
rect 65 840 85 860
rect 105 840 125 860
rect 145 840 165 860
rect 185 840 205 860
rect 225 840 245 860
rect 265 840 285 860
rect 305 840 325 860
rect 345 840 365 860
rect 385 840 405 860
rect 425 840 445 860
rect 465 840 485 860
rect 505 840 525 860
rect 545 840 565 860
rect 585 840 605 860
rect 625 840 645 860
rect 665 840 685 860
rect 705 840 725 860
rect 745 840 765 860
rect 785 840 805 860
rect 850 840 865 860
rect -185 830 865 840
rect -185 790 865 800
rect -185 770 -170 790
rect -135 770 -115 790
rect -95 770 -75 790
rect -55 770 -35 790
rect -15 770 5 790
rect 25 770 45 790
rect 65 770 85 790
rect 105 770 125 790
rect 145 770 165 790
rect 185 770 205 790
rect 225 770 245 790
rect 265 770 285 790
rect 305 770 325 790
rect 345 770 365 790
rect 385 770 405 790
rect 425 770 445 790
rect 465 770 485 790
rect 505 770 525 790
rect 545 770 565 790
rect 585 770 605 790
rect 625 770 645 790
rect 665 770 685 790
rect 705 770 725 790
rect 745 770 765 790
rect 785 770 805 790
rect 850 770 865 790
rect -185 760 865 770
rect -185 720 865 730
rect -185 700 -170 720
rect -135 700 -115 720
rect -95 700 -75 720
rect -55 700 -35 720
rect -15 700 5 720
rect 25 700 45 720
rect 65 700 85 720
rect 105 700 125 720
rect 145 700 165 720
rect 185 700 205 720
rect 225 700 245 720
rect 265 700 285 720
rect 305 700 325 720
rect 345 700 365 720
rect 385 700 405 720
rect 425 700 445 720
rect 465 700 485 720
rect 505 700 525 720
rect 545 700 565 720
rect 585 700 605 720
rect 625 700 645 720
rect 665 700 685 720
rect 705 700 725 720
rect 745 700 765 720
rect 785 700 805 720
rect 850 700 865 720
rect -185 690 865 700
rect -185 650 865 660
rect -185 630 -170 650
rect -135 630 -115 650
rect -95 630 -75 650
rect -55 630 -35 650
rect -15 630 5 650
rect 25 630 45 650
rect 65 630 85 650
rect 105 630 125 650
rect 145 630 165 650
rect 185 630 205 650
rect 225 630 245 650
rect 265 630 285 650
rect 305 630 325 650
rect 345 630 365 650
rect 385 630 405 650
rect 425 630 445 650
rect 465 630 485 650
rect 505 630 525 650
rect 545 630 565 650
rect 585 630 605 650
rect 625 630 645 650
rect 665 630 685 650
rect 705 630 725 650
rect 745 630 765 650
rect 785 630 805 650
rect 850 630 865 650
rect -185 620 865 630
rect -185 580 865 590
rect -185 560 -170 580
rect -135 560 -115 580
rect -95 560 -75 580
rect -55 560 -35 580
rect -15 560 5 580
rect 25 560 45 580
rect 65 560 85 580
rect 105 560 125 580
rect 145 560 165 580
rect 185 560 205 580
rect 225 560 245 580
rect 265 560 285 580
rect 305 560 325 580
rect 345 560 365 580
rect 385 560 405 580
rect 425 560 445 580
rect 465 560 485 580
rect 505 560 525 580
rect 545 560 565 580
rect 585 560 605 580
rect 625 560 645 580
rect 665 560 685 580
rect 705 560 725 580
rect 745 560 765 580
rect 785 560 805 580
rect 850 560 865 580
rect -185 550 865 560
rect 15 485 1015 495
rect 15 465 30 485
rect 65 465 85 485
rect 105 465 125 485
rect 145 465 165 485
rect 185 465 205 485
rect 225 465 245 485
rect 265 465 285 485
rect 305 465 325 485
rect 345 465 365 485
rect 385 465 405 485
rect 425 465 445 485
rect 465 465 485 485
rect 505 465 525 485
rect 545 465 565 485
rect 585 465 605 485
rect 625 465 645 485
rect 665 465 685 485
rect 705 465 725 485
rect 745 465 765 485
rect 785 465 805 485
rect 825 465 845 485
rect 865 465 885 485
rect 905 465 925 485
rect 945 465 965 485
rect 1000 465 1015 485
rect 15 455 1015 465
rect 1035 450 1190 460
rect 1060 430 1080 450
rect 1100 430 1120 450
rect 1140 430 1160 450
rect 1180 430 1190 450
rect 15 415 1015 425
rect 1035 420 1190 430
rect 15 395 30 415
rect 65 395 85 415
rect 105 395 125 415
rect 145 395 165 415
rect 185 395 205 415
rect 225 395 245 415
rect 265 395 285 415
rect 305 395 325 415
rect 345 395 365 415
rect 385 395 405 415
rect 425 395 445 415
rect 465 395 485 415
rect 505 395 525 415
rect 545 395 565 415
rect 585 395 605 415
rect 625 395 645 415
rect 665 395 685 415
rect 705 395 725 415
rect 745 395 765 415
rect 785 395 805 415
rect 825 395 845 415
rect 865 395 885 415
rect 905 395 925 415
rect 945 395 965 415
rect 1000 395 1015 415
rect 15 385 1015 395
rect 1035 380 1190 390
rect 1060 360 1080 380
rect 1100 360 1120 380
rect 1140 360 1160 380
rect 1180 360 1190 380
rect 15 345 1015 355
rect 1035 350 1190 360
rect 15 325 30 345
rect 65 325 85 345
rect 105 325 125 345
rect 145 325 165 345
rect 185 325 205 345
rect 225 325 245 345
rect 265 325 285 345
rect 305 325 325 345
rect 345 325 365 345
rect 385 325 405 345
rect 425 325 445 345
rect 465 325 485 345
rect 505 325 525 345
rect 545 325 565 345
rect 585 325 605 345
rect 625 325 645 345
rect 665 325 685 345
rect 705 325 725 345
rect 745 325 765 345
rect 785 325 805 345
rect 825 325 845 345
rect 865 325 885 345
rect 905 325 925 345
rect 945 325 965 345
rect 1000 325 1015 345
rect 15 315 1015 325
rect 1035 310 1190 320
rect 1060 290 1080 310
rect 1100 290 1120 310
rect 1140 290 1160 310
rect 1180 290 1190 310
rect 15 275 1015 285
rect 1035 280 1190 290
rect 15 255 30 275
rect 65 255 85 275
rect 105 255 125 275
rect 145 255 165 275
rect 185 255 205 275
rect 225 255 245 275
rect 265 255 285 275
rect 305 255 325 275
rect 345 255 365 275
rect 385 255 405 275
rect 425 255 445 275
rect 465 255 485 275
rect 505 255 525 275
rect 545 255 565 275
rect 585 255 605 275
rect 625 255 645 275
rect 665 255 685 275
rect 705 255 725 275
rect 745 255 765 275
rect 785 255 805 275
rect 825 255 845 275
rect 865 255 885 275
rect 905 255 925 275
rect 945 255 965 275
rect 1000 255 1015 275
rect 15 245 1015 255
rect 1035 240 1190 250
rect 1060 220 1080 240
rect 1100 220 1120 240
rect 1140 220 1160 240
rect 1180 220 1190 240
rect 15 205 1015 215
rect 1035 210 1190 220
rect 15 185 30 205
rect 65 185 85 205
rect 105 185 125 205
rect 145 185 165 205
rect 185 185 205 205
rect 225 185 245 205
rect 265 185 285 205
rect 305 185 325 205
rect 345 185 365 205
rect 385 185 405 205
rect 425 185 445 205
rect 465 185 485 205
rect 505 185 525 205
rect 545 185 565 205
rect 585 185 605 205
rect 625 185 645 205
rect 665 185 685 205
rect 705 185 725 205
rect 745 185 765 205
rect 785 185 805 205
rect 825 185 845 205
rect 865 185 885 205
rect 905 185 925 205
rect 945 185 965 205
rect 1000 185 1015 205
rect 15 175 1015 185
rect 1035 170 1190 180
rect 1060 150 1080 170
rect 1100 150 1120 170
rect 1140 150 1160 170
rect 1180 150 1190 170
rect 15 135 1015 145
rect 1035 140 1190 150
rect 15 115 30 135
rect 65 115 85 135
rect 105 115 125 135
rect 145 115 165 135
rect 185 115 205 135
rect 225 115 245 135
rect 265 115 285 135
rect 305 115 325 135
rect 345 115 365 135
rect 385 115 405 135
rect 425 115 445 135
rect 465 115 485 135
rect 505 115 525 135
rect 545 115 565 135
rect 585 115 605 135
rect 625 115 645 135
rect 665 115 685 135
rect 705 115 725 135
rect 745 115 765 135
rect 785 115 805 135
rect 825 115 845 135
rect 865 115 885 135
rect 905 115 925 135
rect 945 115 965 135
rect 1000 115 1015 135
rect 15 105 1015 115
rect 1035 100 1190 110
rect 1060 80 1080 100
rect 1100 80 1120 100
rect 1140 80 1160 100
rect 1180 80 1190 100
rect 15 65 1015 75
rect 1035 70 1190 80
rect 15 45 30 65
rect 65 45 85 65
rect 105 45 125 65
rect 145 45 165 65
rect 185 45 205 65
rect 225 45 245 65
rect 265 45 285 65
rect 305 45 325 65
rect 345 45 365 65
rect 385 45 405 65
rect 425 45 445 65
rect 465 45 485 65
rect 505 45 525 65
rect 545 45 565 65
rect 585 45 605 65
rect 625 45 645 65
rect 665 45 685 65
rect 705 45 725 65
rect 745 45 765 65
rect 785 45 805 65
rect 825 45 845 65
rect 865 45 885 65
rect 905 45 925 65
rect 945 45 965 65
rect 1000 45 1015 65
rect 15 35 1015 45
rect 1035 30 1190 40
rect 1060 10 1080 30
rect 1100 10 1120 30
rect 1140 10 1160 30
rect 1180 10 1190 30
rect 15 -5 1015 5
rect 1035 0 1190 10
rect 15 -25 30 -5
rect 65 -25 85 -5
rect 105 -25 125 -5
rect 145 -25 165 -5
rect 185 -25 205 -5
rect 225 -25 245 -5
rect 265 -25 285 -5
rect 305 -25 325 -5
rect 345 -25 365 -5
rect 385 -25 405 -5
rect 425 -25 445 -5
rect 465 -25 485 -5
rect 505 -25 525 -5
rect 545 -25 565 -5
rect 585 -25 605 -5
rect 625 -25 645 -5
rect 665 -25 685 -5
rect 705 -25 725 -5
rect 745 -25 765 -5
rect 785 -25 805 -5
rect 825 -25 845 -5
rect 865 -25 885 -5
rect 905 -25 925 -5
rect 945 -25 965 -5
rect 1000 -25 1015 -5
rect 15 -35 1015 -25
rect 1035 -40 1190 -30
rect 1060 -60 1080 -40
rect 1100 -60 1120 -40
rect 1140 -60 1160 -40
rect 1180 -60 1190 -40
rect 15 -75 1015 -65
rect 1035 -70 1190 -60
rect 15 -95 30 -75
rect 65 -95 85 -75
rect 105 -95 125 -75
rect 145 -95 165 -75
rect 185 -95 205 -75
rect 225 -95 245 -75
rect 265 -95 285 -75
rect 305 -95 325 -75
rect 345 -95 365 -75
rect 385 -95 405 -75
rect 425 -95 445 -75
rect 465 -95 485 -75
rect 505 -95 525 -75
rect 545 -95 565 -75
rect 585 -95 605 -75
rect 625 -95 645 -75
rect 665 -95 685 -75
rect 705 -95 725 -75
rect 745 -95 765 -75
rect 785 -95 805 -75
rect 825 -95 845 -75
rect 865 -95 885 -75
rect 905 -95 925 -75
rect 945 -95 965 -75
rect 1000 -95 1015 -75
rect 15 -105 1015 -95
rect 1035 -110 1190 -100
rect 1060 -130 1080 -110
rect 1100 -130 1120 -110
rect 1140 -130 1160 -110
rect 1180 -130 1190 -110
rect 15 -145 1015 -135
rect 1035 -140 1190 -130
rect 15 -165 30 -145
rect 65 -165 85 -145
rect 105 -165 125 -145
rect 145 -165 165 -145
rect 185 -165 205 -145
rect 225 -165 245 -145
rect 265 -165 285 -145
rect 305 -165 325 -145
rect 345 -165 365 -145
rect 385 -165 405 -145
rect 425 -165 445 -145
rect 465 -165 485 -145
rect 505 -165 525 -145
rect 545 -165 565 -145
rect 585 -165 605 -145
rect 625 -165 645 -145
rect 665 -165 685 -145
rect 705 -165 725 -145
rect 745 -165 765 -145
rect 785 -165 805 -145
rect 825 -165 845 -145
rect 865 -165 885 -145
rect 905 -165 925 -145
rect 945 -165 965 -145
rect 1000 -165 1015 -145
rect 15 -175 1015 -165
rect 1035 -180 1190 -170
rect 1060 -200 1080 -180
rect 1100 -200 1120 -180
rect 1140 -200 1160 -180
rect 1180 -200 1190 -180
rect 15 -215 1015 -205
rect 1035 -210 1190 -200
rect 15 -235 30 -215
rect 65 -235 85 -215
rect 105 -235 125 -215
rect 145 -235 165 -215
rect 185 -235 205 -215
rect 225 -235 245 -215
rect 265 -235 285 -215
rect 305 -235 325 -215
rect 345 -235 365 -215
rect 385 -235 405 -215
rect 425 -235 445 -215
rect 465 -235 485 -215
rect 505 -235 525 -215
rect 545 -235 565 -215
rect 585 -235 605 -215
rect 625 -235 645 -215
rect 665 -235 685 -215
rect 705 -235 725 -215
rect 745 -235 765 -215
rect 785 -235 805 -215
rect 825 -235 845 -215
rect 865 -235 885 -215
rect 905 -235 925 -215
rect 945 -235 965 -215
rect 1000 -235 1015 -215
rect 15 -245 1015 -235
rect 1035 -250 1190 -240
rect 1060 -270 1080 -250
rect 1100 -270 1120 -250
rect 1140 -270 1160 -250
rect 1180 -270 1190 -250
rect 15 -285 1015 -275
rect 1035 -280 1190 -270
rect 15 -305 30 -285
rect 65 -305 85 -285
rect 105 -305 125 -285
rect 145 -305 165 -285
rect 185 -305 205 -285
rect 225 -305 245 -285
rect 265 -305 285 -285
rect 305 -305 325 -285
rect 345 -305 365 -285
rect 385 -305 405 -285
rect 425 -305 445 -285
rect 465 -305 485 -285
rect 505 -305 525 -285
rect 545 -305 565 -285
rect 585 -305 605 -285
rect 625 -305 645 -285
rect 665 -305 685 -285
rect 705 -305 725 -285
rect 745 -305 765 -285
rect 785 -305 805 -285
rect 825 -305 845 -285
rect 865 -305 885 -285
rect 905 -305 925 -285
rect 945 -305 965 -285
rect 1000 -305 1015 -285
rect 15 -315 1015 -305
rect 1035 -320 1190 -310
rect 1060 -340 1080 -320
rect 1100 -340 1120 -320
rect 1140 -340 1160 -320
rect 1180 -340 1190 -320
rect 15 -355 1015 -345
rect 1035 -350 1190 -340
rect 15 -375 30 -355
rect 65 -375 85 -355
rect 105 -375 125 -355
rect 145 -375 165 -355
rect 185 -375 205 -355
rect 225 -375 245 -355
rect 265 -375 285 -355
rect 305 -375 325 -355
rect 345 -375 365 -355
rect 385 -375 405 -355
rect 425 -375 445 -355
rect 465 -375 485 -355
rect 505 -375 525 -355
rect 545 -375 565 -355
rect 585 -375 605 -355
rect 625 -375 645 -355
rect 665 -375 685 -355
rect 705 -375 725 -355
rect 745 -375 765 -355
rect 785 -375 805 -355
rect 825 -375 845 -355
rect 865 -375 885 -355
rect 905 -375 925 -355
rect 945 -375 965 -355
rect 1000 -375 1015 -355
rect 15 -385 1015 -375
rect 1035 -390 1190 -380
rect 1060 -410 1080 -390
rect 1100 -410 1120 -390
rect 1140 -410 1160 -390
rect 1180 -410 1190 -390
rect 15 -425 1015 -415
rect 1035 -420 1190 -410
rect 15 -445 30 -425
rect 65 -445 85 -425
rect 105 -445 125 -425
rect 145 -445 165 -425
rect 185 -445 205 -425
rect 225 -445 245 -425
rect 265 -445 285 -425
rect 305 -445 325 -425
rect 345 -445 365 -425
rect 385 -445 405 -425
rect 425 -445 445 -425
rect 465 -445 485 -425
rect 505 -445 525 -425
rect 545 -445 565 -425
rect 585 -445 605 -425
rect 625 -445 645 -425
rect 665 -445 685 -425
rect 705 -445 725 -425
rect 745 -445 765 -425
rect 785 -445 805 -425
rect 825 -445 845 -425
rect 865 -445 885 -425
rect 905 -445 925 -425
rect 945 -445 965 -425
rect 1000 -445 1015 -425
rect 15 -455 1015 -445
rect 1035 -460 1190 -450
rect 1060 -480 1080 -460
rect 1100 -480 1120 -460
rect 1140 -480 1160 -460
rect 1180 -480 1190 -460
rect 15 -495 1015 -485
rect 1035 -490 1190 -480
rect 15 -515 30 -495
rect 65 -515 85 -495
rect 105 -515 125 -495
rect 145 -515 165 -495
rect 185 -515 205 -495
rect 225 -515 245 -495
rect 265 -515 285 -495
rect 305 -515 325 -495
rect 345 -515 365 -495
rect 385 -515 405 -495
rect 425 -515 445 -495
rect 465 -515 485 -495
rect 505 -515 525 -495
rect 545 -515 565 -495
rect 585 -515 605 -495
rect 625 -515 645 -495
rect 665 -515 685 -495
rect 705 -515 725 -495
rect 745 -515 765 -495
rect 785 -515 805 -495
rect 825 -515 845 -495
rect 865 -515 885 -495
rect 905 -515 925 -495
rect 945 -515 965 -495
rect 1000 -515 1015 -495
rect 15 -525 1015 -515
rect 1035 -530 1190 -520
rect 1060 -550 1080 -530
rect 1100 -550 1120 -530
rect 1140 -550 1160 -530
rect 1180 -550 1190 -530
rect 15 -565 1015 -555
rect 1035 -560 1190 -550
rect 15 -585 30 -565
rect 65 -585 85 -565
rect 105 -585 125 -565
rect 145 -585 165 -565
rect 185 -585 205 -565
rect 225 -585 245 -565
rect 265 -585 285 -565
rect 305 -585 325 -565
rect 345 -585 365 -565
rect 385 -585 405 -565
rect 425 -585 445 -565
rect 465 -585 485 -565
rect 505 -585 525 -565
rect 545 -585 565 -565
rect 585 -585 605 -565
rect 625 -585 645 -565
rect 665 -585 685 -565
rect 705 -585 725 -565
rect 745 -585 765 -565
rect 785 -585 805 -565
rect 825 -585 845 -565
rect 865 -585 885 -565
rect 905 -585 925 -565
rect 945 -585 965 -565
rect 1000 -585 1015 -565
rect 15 -595 1015 -585
rect -135 -635 1165 -625
rect -135 -655 -120 -635
rect -95 -655 -75 -635
rect -55 -655 -35 -635
rect -15 -655 5 -635
rect 25 -655 45 -635
rect 65 -655 85 -635
rect 105 -655 125 -635
rect 145 -655 165 -635
rect 185 -655 205 -635
rect 225 -655 245 -635
rect 265 -655 285 -635
rect 305 -655 325 -635
rect 345 -655 365 -635
rect 385 -655 405 -635
rect 425 -655 445 -635
rect 465 -655 485 -635
rect 505 -655 525 -635
rect 545 -655 565 -635
rect 585 -655 605 -635
rect 625 -655 645 -635
rect 665 -655 685 -635
rect 705 -655 725 -635
rect 745 -655 765 -635
rect 785 -655 805 -635
rect 825 -655 845 -635
rect 865 -655 885 -635
rect 905 -655 925 -635
rect 945 -655 965 -635
rect 985 -655 1005 -635
rect 1025 -655 1045 -635
rect 1065 -655 1085 -635
rect 1105 -655 1125 -635
rect 1150 -655 1165 -635
rect -135 -675 1165 -655
rect -135 -695 -120 -675
rect -95 -695 -75 -675
rect -55 -695 -35 -675
rect -15 -695 5 -675
rect 25 -695 45 -675
rect 65 -695 85 -675
rect 105 -695 125 -675
rect 145 -695 165 -675
rect 185 -695 205 -675
rect 225 -695 245 -675
rect 265 -695 285 -675
rect 305 -695 325 -675
rect 345 -695 365 -675
rect 385 -695 405 -675
rect 425 -695 445 -675
rect 465 -695 485 -675
rect 505 -695 525 -675
rect 545 -695 565 -675
rect 585 -695 605 -675
rect 625 -695 645 -675
rect 665 -695 685 -675
rect 705 -695 725 -675
rect 745 -695 765 -675
rect 785 -695 805 -675
rect 825 -695 845 -675
rect 865 -695 885 -675
rect 905 -695 925 -675
rect 945 -695 965 -675
rect 985 -695 1005 -675
rect 1025 -695 1045 -675
rect 1065 -695 1085 -675
rect 1105 -695 1125 -675
rect 1150 -695 1165 -675
rect -135 -705 1165 -695
rect -310 -720 -155 -710
rect -310 -750 -300 -720
rect -280 -750 -260 -720
rect -240 -750 -220 -720
rect -200 -750 -180 -720
rect -310 -760 -155 -750
rect -135 -775 1165 -765
rect -135 -795 -120 -775
rect -95 -795 -75 -775
rect -55 -795 -35 -775
rect -15 -795 5 -775
rect 25 -795 45 -775
rect 65 -795 85 -775
rect 105 -795 125 -775
rect 145 -795 165 -775
rect 185 -795 205 -775
rect 225 -795 245 -775
rect 265 -795 285 -775
rect 305 -795 325 -775
rect 345 -795 365 -775
rect 385 -795 405 -775
rect 425 -795 445 -775
rect 465 -795 485 -775
rect 505 -795 525 -775
rect 545 -795 565 -775
rect 585 -795 605 -775
rect 625 -795 645 -775
rect 665 -795 685 -775
rect 705 -795 725 -775
rect 745 -795 765 -775
rect 785 -795 805 -775
rect 825 -795 845 -775
rect 865 -795 885 -775
rect 905 -795 925 -775
rect 945 -795 965 -775
rect 985 -795 1005 -775
rect 1025 -795 1045 -775
rect 1065 -795 1085 -775
rect 1105 -795 1125 -775
rect 1150 -795 1165 -775
rect -135 -805 1165 -795
rect -310 -820 -155 -810
rect -310 -850 -300 -820
rect -280 -850 -260 -820
rect -240 -850 -220 -820
rect -200 -850 -180 -820
rect -310 -860 -155 -850
rect -135 -875 1165 -865
rect -135 -895 -120 -875
rect -95 -895 -75 -875
rect -55 -895 -35 -875
rect -15 -895 5 -875
rect 25 -895 45 -875
rect 65 -895 85 -875
rect 105 -895 125 -875
rect 145 -895 165 -875
rect 185 -895 205 -875
rect 225 -895 245 -875
rect 265 -895 285 -875
rect 305 -895 325 -875
rect 345 -895 365 -875
rect 385 -895 405 -875
rect 425 -895 445 -875
rect 465 -895 485 -875
rect 505 -895 525 -875
rect 545 -895 565 -875
rect 585 -895 605 -875
rect 625 -895 645 -875
rect 665 -895 685 -875
rect 705 -895 725 -875
rect 745 -895 765 -875
rect 785 -895 805 -875
rect 825 -895 845 -875
rect 865 -895 885 -875
rect 905 -895 925 -875
rect 945 -895 965 -875
rect 985 -895 1005 -875
rect 1025 -895 1045 -875
rect 1065 -895 1085 -875
rect 1105 -895 1125 -875
rect 1150 -895 1165 -875
rect -135 -905 1165 -895
rect -310 -920 -155 -910
rect -310 -950 -300 -920
rect -280 -950 -260 -920
rect -240 -950 -220 -920
rect -200 -950 -180 -920
rect -310 -960 -155 -950
rect -135 -975 1165 -965
rect -135 -995 -120 -975
rect -95 -995 -75 -975
rect -55 -995 -35 -975
rect -15 -995 5 -975
rect 25 -995 45 -975
rect 65 -995 85 -975
rect 105 -995 125 -975
rect 145 -995 165 -975
rect 185 -995 205 -975
rect 225 -995 245 -975
rect 265 -995 285 -975
rect 305 -995 325 -975
rect 345 -995 365 -975
rect 385 -995 405 -975
rect 425 -995 445 -975
rect 465 -995 485 -975
rect 505 -995 525 -975
rect 545 -995 565 -975
rect 585 -995 605 -975
rect 625 -995 645 -975
rect 665 -995 685 -975
rect 705 -995 725 -975
rect 745 -995 765 -975
rect 785 -995 805 -975
rect 825 -995 845 -975
rect 865 -995 885 -975
rect 905 -995 925 -975
rect 945 -995 965 -975
rect 985 -995 1005 -975
rect 1025 -995 1045 -975
rect 1065 -995 1085 -975
rect 1105 -995 1125 -975
rect 1150 -995 1165 -975
rect -135 -1005 1165 -995
rect -310 -1020 -155 -1010
rect -310 -1050 -300 -1020
rect -280 -1050 -260 -1020
rect -240 -1050 -220 -1020
rect -200 -1050 -180 -1020
rect -310 -1060 -155 -1050
rect -135 -1075 1165 -1065
rect -135 -1095 -120 -1075
rect -95 -1095 -75 -1075
rect -55 -1095 -35 -1075
rect -15 -1095 5 -1075
rect 25 -1095 45 -1075
rect 65 -1095 85 -1075
rect 105 -1095 125 -1075
rect 145 -1095 165 -1075
rect 185 -1095 205 -1075
rect 225 -1095 245 -1075
rect 265 -1095 285 -1075
rect 305 -1095 325 -1075
rect 345 -1095 365 -1075
rect 385 -1095 405 -1075
rect 425 -1095 445 -1075
rect 465 -1095 485 -1075
rect 505 -1095 525 -1075
rect 545 -1095 565 -1075
rect 585 -1095 605 -1075
rect 625 -1095 645 -1075
rect 665 -1095 685 -1075
rect 705 -1095 725 -1075
rect 745 -1095 765 -1075
rect 785 -1095 805 -1075
rect 825 -1095 845 -1075
rect 865 -1095 885 -1075
rect 905 -1095 925 -1075
rect 945 -1095 965 -1075
rect 985 -1095 1005 -1075
rect 1025 -1095 1045 -1075
rect 1065 -1095 1085 -1075
rect 1105 -1095 1125 -1075
rect 1150 -1095 1165 -1075
rect -135 -1105 1165 -1095
rect -310 -1120 -155 -1110
rect -310 -1150 -300 -1120
rect -280 -1150 -260 -1120
rect -240 -1150 -220 -1120
rect -200 -1150 -180 -1120
rect -310 -1160 -155 -1150
rect -135 -1175 1165 -1165
rect -135 -1195 -120 -1175
rect -95 -1195 -75 -1175
rect -55 -1195 -35 -1175
rect -15 -1195 5 -1175
rect 25 -1195 45 -1175
rect 65 -1195 85 -1175
rect 105 -1195 125 -1175
rect 145 -1195 165 -1175
rect 185 -1195 205 -1175
rect 225 -1195 245 -1175
rect 265 -1195 285 -1175
rect 305 -1195 325 -1175
rect 345 -1195 365 -1175
rect 385 -1195 405 -1175
rect 425 -1195 445 -1175
rect 465 -1195 485 -1175
rect 505 -1195 525 -1175
rect 545 -1195 565 -1175
rect 585 -1195 605 -1175
rect 625 -1195 645 -1175
rect 665 -1195 685 -1175
rect 705 -1195 725 -1175
rect 745 -1195 765 -1175
rect 785 -1195 805 -1175
rect 825 -1195 845 -1175
rect 865 -1195 885 -1175
rect 905 -1195 925 -1175
rect 945 -1195 965 -1175
rect 985 -1195 1005 -1175
rect 1025 -1195 1045 -1175
rect 1065 -1195 1085 -1175
rect 1105 -1195 1125 -1175
rect 1150 -1195 1165 -1175
rect -135 -1205 1165 -1195
<< viali >>
rect 125 880 145 900
rect 165 880 185 900
rect 205 880 225 900
rect 245 880 265 900
rect 285 880 305 900
rect 325 880 345 900
rect 485 770 505 790
rect 525 770 545 790
rect 565 770 585 790
rect 605 770 625 790
rect 645 770 665 790
rect 685 770 705 790
rect 125 700 145 720
rect 165 700 185 720
rect 205 700 225 720
rect 245 700 265 720
rect 285 700 305 720
rect 325 700 345 720
rect 485 630 505 650
rect 525 630 545 650
rect 565 630 585 650
rect 605 630 625 650
rect 645 630 665 650
rect 685 630 705 650
rect 125 560 145 580
rect 165 560 185 580
rect 205 560 225 580
rect 245 560 265 580
rect 285 560 305 580
rect 325 560 345 580
rect 165 465 185 485
rect 205 465 225 485
rect 245 465 265 485
rect 285 465 305 485
rect 325 465 345 485
rect 365 465 385 485
rect 1040 430 1060 450
rect 1080 430 1100 450
rect 1120 430 1140 450
rect 1160 430 1180 450
rect 485 395 505 415
rect 525 395 545 415
rect 565 395 585 415
rect 605 395 625 415
rect 645 395 665 415
rect 685 395 705 415
rect 1040 360 1060 380
rect 1080 360 1100 380
rect 1120 360 1140 380
rect 1160 360 1180 380
rect 165 325 185 345
rect 205 325 225 345
rect 245 325 265 345
rect 285 325 305 345
rect 325 325 345 345
rect 365 325 385 345
rect 1040 290 1060 310
rect 1080 290 1100 310
rect 1120 290 1140 310
rect 1160 290 1180 310
rect 485 255 505 275
rect 525 255 545 275
rect 565 255 585 275
rect 605 255 625 275
rect 645 255 665 275
rect 685 255 705 275
rect 1040 220 1060 240
rect 1080 220 1100 240
rect 1120 220 1140 240
rect 1160 220 1180 240
rect 165 185 185 205
rect 205 185 225 205
rect 245 185 265 205
rect 285 185 305 205
rect 325 185 345 205
rect 365 185 385 205
rect 1040 150 1060 170
rect 1080 150 1100 170
rect 1120 150 1140 170
rect 1160 150 1180 170
rect 485 115 505 135
rect 525 115 545 135
rect 565 115 585 135
rect 605 115 625 135
rect 645 115 665 135
rect 685 115 705 135
rect 1040 80 1060 100
rect 1080 80 1100 100
rect 1120 80 1140 100
rect 1160 80 1180 100
rect 165 45 185 65
rect 205 45 225 65
rect 245 45 265 65
rect 285 45 305 65
rect 325 45 345 65
rect 365 45 385 65
rect 1040 10 1060 30
rect 1080 10 1100 30
rect 1120 10 1140 30
rect 1160 10 1180 30
rect 485 -25 505 -5
rect 525 -25 545 -5
rect 565 -25 585 -5
rect 605 -25 625 -5
rect 645 -25 665 -5
rect 685 -25 705 -5
rect 1040 -60 1060 -40
rect 1080 -60 1100 -40
rect 1120 -60 1140 -40
rect 1160 -60 1180 -40
rect 165 -95 185 -75
rect 205 -95 225 -75
rect 245 -95 265 -75
rect 285 -95 305 -75
rect 325 -95 345 -75
rect 365 -95 385 -75
rect 1040 -130 1060 -110
rect 1080 -130 1100 -110
rect 1120 -130 1140 -110
rect 1160 -130 1180 -110
rect 485 -165 505 -145
rect 525 -165 545 -145
rect 565 -165 585 -145
rect 605 -165 625 -145
rect 645 -165 665 -145
rect 685 -165 705 -145
rect 1040 -200 1060 -180
rect 1080 -200 1100 -180
rect 1120 -200 1140 -180
rect 1160 -200 1180 -180
rect 165 -235 185 -215
rect 205 -235 225 -215
rect 245 -235 265 -215
rect 285 -235 305 -215
rect 325 -235 345 -215
rect 365 -235 385 -215
rect 1040 -270 1060 -250
rect 1080 -270 1100 -250
rect 1120 -270 1140 -250
rect 1160 -270 1180 -250
rect 485 -305 505 -285
rect 525 -305 545 -285
rect 565 -305 585 -285
rect 605 -305 625 -285
rect 645 -305 665 -285
rect 685 -305 705 -285
rect 1040 -340 1060 -320
rect 1080 -340 1100 -320
rect 1120 -340 1140 -320
rect 1160 -340 1180 -320
rect 165 -375 185 -355
rect 205 -375 225 -355
rect 245 -375 265 -355
rect 285 -375 305 -355
rect 325 -375 345 -355
rect 365 -375 385 -355
rect 1040 -410 1060 -390
rect 1080 -410 1100 -390
rect 1120 -410 1140 -390
rect 1160 -410 1180 -390
rect 485 -445 505 -425
rect 525 -445 545 -425
rect 565 -445 585 -425
rect 605 -445 625 -425
rect 645 -445 665 -425
rect 685 -445 705 -425
rect 1040 -480 1060 -460
rect 1080 -480 1100 -460
rect 1120 -480 1140 -460
rect 1160 -480 1180 -460
rect 165 -515 185 -495
rect 205 -515 225 -495
rect 245 -515 265 -495
rect 285 -515 305 -495
rect 325 -515 345 -495
rect 365 -515 385 -495
rect 1040 -550 1060 -530
rect 1080 -550 1100 -530
rect 1120 -550 1140 -530
rect 1160 -550 1180 -530
rect 485 -585 505 -565
rect 525 -585 545 -565
rect 565 -585 585 -565
rect 605 -585 625 -565
rect 645 -585 665 -565
rect 685 -585 705 -565
rect 645 -655 665 -635
rect 685 -655 705 -635
rect 725 -655 745 -635
rect 765 -655 785 -635
rect 805 -655 825 -635
rect 845 -655 865 -635
rect 645 -695 665 -675
rect 685 -695 705 -675
rect 725 -695 745 -675
rect 765 -695 785 -675
rect 805 -695 825 -675
rect 845 -695 865 -675
rect -300 -750 -280 -720
rect -260 -750 -240 -720
rect -220 -750 -200 -720
rect -180 -750 -160 -720
rect 165 -795 185 -775
rect 205 -795 225 -775
rect 245 -795 265 -775
rect 285 -795 305 -775
rect 325 -795 345 -775
rect 365 -795 385 -775
rect -300 -850 -280 -820
rect -260 -850 -240 -820
rect -220 -850 -200 -820
rect -180 -850 -160 -820
rect 645 -895 665 -875
rect 685 -895 705 -875
rect 725 -895 745 -875
rect 765 -895 785 -875
rect 805 -895 825 -875
rect 845 -895 865 -875
rect -300 -950 -280 -920
rect -260 -950 -240 -920
rect -220 -950 -200 -920
rect -180 -950 -160 -920
rect 165 -995 185 -975
rect 205 -995 225 -975
rect 245 -995 265 -975
rect 285 -995 305 -975
rect 325 -995 345 -975
rect 365 -995 385 -975
rect -300 -1050 -280 -1020
rect -260 -1050 -240 -1020
rect -220 -1050 -200 -1020
rect -180 -1050 -160 -1020
rect 645 -1095 665 -1075
rect 685 -1095 705 -1075
rect 725 -1095 745 -1075
rect 765 -1095 785 -1075
rect 805 -1095 825 -1075
rect 845 -1095 865 -1075
rect -300 -1150 -280 -1120
rect -260 -1150 -240 -1120
rect -220 -1150 -200 -1120
rect -180 -1150 -160 -1120
rect 165 -1195 185 -1175
rect 205 -1195 225 -1175
rect 245 -1195 265 -1175
rect 285 -1195 305 -1175
rect 325 -1195 345 -1175
rect 365 -1195 385 -1175
<< metal1 >>
rect 115 900 355 925
rect 115 880 125 900
rect 145 880 165 900
rect 185 880 205 900
rect 225 880 245 900
rect 265 880 285 900
rect 305 880 325 900
rect 345 880 355 900
rect 115 720 355 880
rect 115 700 125 720
rect 145 700 165 720
rect 185 700 205 720
rect 225 700 245 720
rect 265 700 285 720
rect 305 700 325 720
rect 345 700 355 720
rect 115 580 355 700
rect 115 560 125 580
rect 145 560 165 580
rect 185 560 205 580
rect 225 560 245 580
rect 265 560 285 580
rect 305 560 325 580
rect 345 560 355 580
rect 115 550 355 560
rect 475 790 715 800
rect 475 770 485 790
rect 505 770 525 790
rect 545 770 565 790
rect 585 770 605 790
rect 625 770 645 790
rect 665 770 685 790
rect 705 770 715 790
rect 475 650 715 770
rect 475 630 485 650
rect 505 630 525 650
rect 545 630 565 650
rect 585 630 605 650
rect 625 630 645 650
rect 665 630 685 650
rect 705 630 715 650
rect 155 485 395 495
rect 155 465 165 485
rect 185 465 205 485
rect 225 465 245 485
rect 265 465 285 485
rect 305 465 325 485
rect 345 465 365 485
rect 385 465 395 485
rect 155 345 395 465
rect 155 325 165 345
rect 185 325 205 345
rect 225 325 245 345
rect 265 325 285 345
rect 305 325 325 345
rect 345 325 365 345
rect 385 325 395 345
rect 155 205 395 325
rect 155 185 165 205
rect 185 185 205 205
rect 225 185 245 205
rect 265 185 285 205
rect 305 185 325 205
rect 345 185 365 205
rect 385 185 395 205
rect 155 65 395 185
rect 155 45 165 65
rect 185 45 205 65
rect 225 45 245 65
rect 265 45 285 65
rect 305 45 325 65
rect 345 45 365 65
rect 385 45 395 65
rect 155 -75 395 45
rect 155 -95 165 -75
rect 185 -95 205 -75
rect 225 -95 245 -75
rect 265 -95 285 -75
rect 305 -95 325 -75
rect 345 -95 365 -75
rect 385 -95 395 -75
rect 155 -215 395 -95
rect 155 -235 165 -215
rect 185 -235 205 -215
rect 225 -235 245 -215
rect 265 -235 285 -215
rect 305 -235 325 -215
rect 345 -235 365 -215
rect 385 -235 395 -215
rect 155 -355 395 -235
rect 155 -375 165 -355
rect 185 -375 205 -355
rect 225 -375 245 -355
rect 265 -375 285 -355
rect 305 -375 325 -355
rect 345 -375 365 -355
rect 385 -375 395 -355
rect 155 -495 395 -375
rect 155 -515 165 -495
rect 185 -515 205 -495
rect 225 -515 245 -495
rect 265 -515 285 -495
rect 305 -515 325 -495
rect 345 -515 365 -495
rect 385 -515 395 -495
rect -310 -720 -145 -710
rect -310 -750 -300 -720
rect -280 -750 -260 -720
rect -240 -750 -220 -720
rect -200 -750 -180 -720
rect -160 -750 -145 -720
rect -310 -820 -145 -750
rect -310 -850 -300 -820
rect -280 -850 -260 -820
rect -240 -850 -220 -820
rect -200 -850 -180 -820
rect -160 -850 -145 -820
rect -310 -920 -145 -850
rect -310 -950 -300 -920
rect -280 -950 -260 -920
rect -240 -950 -220 -920
rect -200 -950 -180 -920
rect -160 -950 -145 -920
rect -310 -1020 -145 -950
rect -310 -1050 -300 -1020
rect -280 -1050 -260 -1020
rect -240 -1050 -220 -1020
rect -200 -1050 -180 -1020
rect -160 -1050 -145 -1020
rect -310 -1120 -145 -1050
rect -310 -1150 -300 -1120
rect -280 -1150 -260 -1120
rect -240 -1150 -220 -1120
rect -200 -1150 -180 -1120
rect -160 -1150 -145 -1120
rect -310 -1160 -145 -1150
rect 155 -775 395 -515
rect 475 415 715 630
rect 475 395 485 415
rect 505 395 525 415
rect 545 395 565 415
rect 585 395 605 415
rect 625 395 645 415
rect 665 395 685 415
rect 705 395 715 415
rect 475 275 715 395
rect 475 255 485 275
rect 505 255 525 275
rect 545 255 565 275
rect 585 255 605 275
rect 625 255 645 275
rect 665 255 685 275
rect 705 255 715 275
rect 475 135 715 255
rect 475 115 485 135
rect 505 115 525 135
rect 545 115 565 135
rect 585 115 605 135
rect 625 115 645 135
rect 665 115 685 135
rect 705 115 715 135
rect 475 -5 715 115
rect 475 -25 485 -5
rect 505 -25 525 -5
rect 545 -25 565 -5
rect 585 -25 605 -5
rect 625 -25 645 -5
rect 665 -25 685 -5
rect 705 -25 715 -5
rect 475 -145 715 -25
rect 475 -165 485 -145
rect 505 -165 525 -145
rect 545 -165 565 -145
rect 585 -165 605 -145
rect 625 -165 645 -145
rect 665 -165 685 -145
rect 705 -165 715 -145
rect 475 -285 715 -165
rect 475 -305 485 -285
rect 505 -305 525 -285
rect 545 -305 565 -285
rect 585 -305 605 -285
rect 625 -305 645 -285
rect 665 -305 685 -285
rect 705 -305 715 -285
rect 475 -425 715 -305
rect 475 -445 485 -425
rect 505 -445 525 -425
rect 545 -445 565 -425
rect 585 -445 605 -425
rect 625 -445 645 -425
rect 665 -445 685 -425
rect 705 -445 715 -425
rect 475 -565 715 -445
rect 1025 450 1190 460
rect 1025 430 1040 450
rect 1060 430 1080 450
rect 1100 430 1120 450
rect 1140 430 1160 450
rect 1180 430 1190 450
rect 1025 380 1190 430
rect 1025 360 1040 380
rect 1060 360 1080 380
rect 1100 360 1120 380
rect 1140 360 1160 380
rect 1180 360 1190 380
rect 1025 310 1190 360
rect 1025 290 1040 310
rect 1060 290 1080 310
rect 1100 290 1120 310
rect 1140 290 1160 310
rect 1180 290 1190 310
rect 1025 240 1190 290
rect 1025 220 1040 240
rect 1060 220 1080 240
rect 1100 220 1120 240
rect 1140 220 1160 240
rect 1180 220 1190 240
rect 1025 170 1190 220
rect 1025 150 1040 170
rect 1060 150 1080 170
rect 1100 150 1120 170
rect 1140 150 1160 170
rect 1180 150 1190 170
rect 1025 100 1190 150
rect 1025 80 1040 100
rect 1060 80 1080 100
rect 1100 80 1120 100
rect 1140 80 1160 100
rect 1180 80 1190 100
rect 1025 30 1190 80
rect 1025 10 1040 30
rect 1060 10 1080 30
rect 1100 10 1120 30
rect 1140 10 1160 30
rect 1180 10 1190 30
rect 1025 -40 1190 10
rect 1025 -60 1040 -40
rect 1060 -60 1080 -40
rect 1100 -60 1120 -40
rect 1140 -60 1160 -40
rect 1180 -60 1190 -40
rect 1025 -110 1190 -60
rect 1025 -130 1040 -110
rect 1060 -130 1080 -110
rect 1100 -130 1120 -110
rect 1140 -130 1160 -110
rect 1180 -130 1190 -110
rect 1025 -180 1190 -130
rect 1025 -200 1040 -180
rect 1060 -200 1080 -180
rect 1100 -200 1120 -180
rect 1140 -200 1160 -180
rect 1180 -200 1190 -180
rect 1025 -250 1190 -200
rect 1025 -270 1040 -250
rect 1060 -270 1080 -250
rect 1100 -270 1120 -250
rect 1140 -270 1160 -250
rect 1180 -270 1190 -250
rect 1025 -320 1190 -270
rect 1025 -340 1040 -320
rect 1060 -340 1080 -320
rect 1100 -340 1120 -320
rect 1140 -340 1160 -320
rect 1180 -340 1190 -320
rect 1025 -390 1190 -340
rect 1025 -410 1040 -390
rect 1060 -410 1080 -390
rect 1100 -410 1120 -390
rect 1140 -410 1160 -390
rect 1180 -410 1190 -390
rect 1025 -460 1190 -410
rect 1025 -480 1040 -460
rect 1060 -480 1080 -460
rect 1100 -480 1120 -460
rect 1140 -480 1160 -460
rect 1180 -480 1190 -460
rect 1025 -530 1190 -480
rect 1025 -550 1040 -530
rect 1060 -550 1080 -530
rect 1100 -550 1120 -530
rect 1140 -550 1160 -530
rect 1180 -550 1190 -530
rect 1025 -560 1190 -550
rect 475 -585 485 -565
rect 505 -585 525 -565
rect 545 -585 565 -565
rect 585 -585 605 -565
rect 625 -585 645 -565
rect 665 -585 685 -565
rect 705 -585 715 -565
rect 475 -595 715 -585
rect 155 -795 165 -775
rect 185 -795 205 -775
rect 225 -795 245 -775
rect 265 -795 285 -775
rect 305 -795 325 -775
rect 345 -795 365 -775
rect 385 -795 395 -775
rect 155 -975 395 -795
rect 155 -995 165 -975
rect 185 -995 205 -975
rect 225 -995 245 -975
rect 265 -995 285 -975
rect 305 -995 325 -975
rect 345 -995 365 -975
rect 385 -995 395 -975
rect 155 -1175 395 -995
rect 155 -1195 165 -1175
rect 185 -1195 205 -1175
rect 225 -1195 245 -1175
rect 265 -1195 285 -1175
rect 305 -1195 325 -1175
rect 345 -1195 365 -1175
rect 385 -1195 395 -1175
rect 155 -1205 395 -1195
rect 635 -635 875 -625
rect 635 -655 645 -635
rect 665 -655 685 -635
rect 705 -655 725 -635
rect 745 -655 765 -635
rect 785 -655 805 -635
rect 825 -655 845 -635
rect 865 -655 875 -635
rect 635 -675 875 -655
rect 635 -695 645 -675
rect 665 -695 685 -675
rect 705 -695 725 -675
rect 745 -695 765 -675
rect 785 -695 805 -675
rect 825 -695 845 -675
rect 865 -695 875 -675
rect 635 -875 875 -695
rect 635 -895 645 -875
rect 665 -895 685 -875
rect 705 -895 725 -875
rect 745 -895 765 -875
rect 785 -895 805 -875
rect 825 -895 845 -875
rect 865 -895 875 -875
rect 635 -1075 875 -895
rect 635 -1095 645 -1075
rect 665 -1095 685 -1075
rect 705 -1095 725 -1075
rect 745 -1095 765 -1075
rect 785 -1095 805 -1075
rect 825 -1095 845 -1075
rect 865 -1095 875 -1075
rect 635 -1220 875 -1095
<< labels >>
rlabel metal1 755 -1215 755 -1215 1 GND
port 7 n
rlabel metal1 260 -605 260 -605 1 res
port 9 n
rlabel metal1 1185 -50 1185 -50 1 Vin
port 11 n
rlabel metal1 -305 -935 -305 -935 1 Vb3
port 10 n
rlabel metal1 210 915 210 915 1 VDD
port 2 n
rlabel metal1 590 520 590 520 1 Vout
port 8 n
rlabel poly -210 715 -210 715 1 diode
port 12 n
<< end >>
