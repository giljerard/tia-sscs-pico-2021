magic
tech sky130A
timestamp 1634683452
<< xpolycontact >>
rect -1480 1174 -1240 1315
rect -1099 1174 -860 1315
<< xpolyres >>
rect -1240 1174 -1099 1315
<< viali >>
rect -1470 1274 -1450 1294
rect -1430 1274 -1410 1294
rect -1390 1274 -1370 1294
rect -1350 1274 -1330 1294
rect -1310 1274 -1290 1294
rect -1270 1274 -1250 1294
rect -1470 1234 -1450 1254
rect -1430 1234 -1410 1254
rect -1390 1234 -1370 1254
rect -1350 1234 -1330 1254
rect -1310 1234 -1290 1254
rect -1270 1234 -1250 1254
rect -1470 1194 -1450 1214
rect -1430 1194 -1410 1214
rect -1390 1194 -1370 1214
rect -1350 1194 -1330 1214
rect -1310 1194 -1290 1214
rect -1270 1194 -1250 1214
rect -1090 1274 -1070 1294
rect -1050 1274 -1030 1294
rect -1010 1274 -990 1294
rect -970 1274 -950 1294
rect -930 1274 -910 1294
rect -890 1274 -870 1294
rect -1090 1234 -1070 1254
rect -1050 1234 -1030 1254
rect -1010 1234 -990 1254
rect -970 1234 -950 1254
rect -930 1234 -910 1254
rect -890 1234 -870 1254
rect -1090 1194 -1070 1214
rect -1050 1194 -1030 1214
rect -1010 1194 -990 1214
rect -970 1194 -950 1214
rect -930 1194 -910 1214
rect -890 1194 -870 1214
<< metal1 >>
rect -1480 1294 -1240 1315
rect -1480 1234 -1470 1294
rect -1450 1275 -1430 1294
rect -1410 1275 -1390 1294
rect -1370 1275 -1350 1294
rect -1330 1275 -1310 1294
rect -1290 1275 -1270 1294
rect -1435 1274 -1430 1275
rect -1370 1274 -1360 1275
rect -1325 1274 -1310 1275
rect -1250 1274 -1240 1294
rect -1435 1254 -1415 1274
rect -1380 1254 -1360 1274
rect -1325 1254 -1305 1274
rect -1270 1254 -1240 1274
rect -1435 1240 -1430 1254
rect -1370 1240 -1360 1254
rect -1325 1240 -1310 1254
rect -1450 1234 -1430 1240
rect -1410 1234 -1390 1240
rect -1370 1234 -1350 1240
rect -1330 1234 -1310 1240
rect -1290 1234 -1270 1240
rect -1250 1234 -1240 1254
rect -1480 1220 -1240 1234
rect -1480 1185 -1470 1220
rect -1435 1214 -1415 1220
rect -1380 1214 -1360 1220
rect -1325 1214 -1305 1220
rect -1270 1214 -1240 1220
rect -1435 1194 -1430 1214
rect -1370 1194 -1360 1214
rect -1325 1194 -1310 1214
rect -1250 1194 -1240 1214
rect -1435 1185 -1415 1194
rect -1380 1185 -1360 1194
rect -1325 1185 -1305 1194
rect -1270 1185 -1240 1194
rect -1480 1174 -1240 1185
rect -1099 1305 -860 1315
rect -1099 1294 -1085 1305
rect -1050 1294 -1030 1305
rect -995 1294 -975 1305
rect -940 1294 -920 1305
rect -885 1294 -860 1305
rect -1099 1274 -1090 1294
rect -990 1274 -975 1294
rect -940 1274 -930 1294
rect -870 1274 -860 1294
rect -1099 1270 -1085 1274
rect -1050 1270 -1030 1274
rect -995 1270 -975 1274
rect -940 1270 -920 1274
rect -885 1270 -860 1274
rect -1099 1254 -860 1270
rect -1099 1234 -1090 1254
rect -1070 1250 -1050 1254
rect -1030 1250 -1010 1254
rect -990 1250 -970 1254
rect -950 1250 -930 1254
rect -910 1250 -890 1254
rect -990 1234 -975 1250
rect -940 1234 -930 1250
rect -870 1234 -860 1254
rect -1099 1215 -1085 1234
rect -1050 1215 -1030 1234
rect -995 1215 -975 1234
rect -940 1215 -920 1234
rect -885 1215 -860 1234
rect -1099 1214 -860 1215
rect -1099 1194 -1090 1214
rect -1070 1194 -1050 1214
rect -1030 1194 -1010 1214
rect -990 1194 -970 1214
rect -950 1194 -930 1214
rect -910 1194 -890 1214
rect -870 1194 -860 1214
rect -1099 1174 -860 1194
<< via1 >>
rect -1470 1274 -1450 1275
rect -1450 1274 -1435 1275
rect -1415 1274 -1410 1275
rect -1410 1274 -1390 1275
rect -1390 1274 -1380 1275
rect -1360 1274 -1350 1275
rect -1350 1274 -1330 1275
rect -1330 1274 -1325 1275
rect -1305 1274 -1290 1275
rect -1290 1274 -1270 1275
rect -1470 1254 -1435 1274
rect -1415 1254 -1380 1274
rect -1360 1254 -1325 1274
rect -1305 1254 -1270 1274
rect -1470 1240 -1450 1254
rect -1450 1240 -1435 1254
rect -1415 1240 -1410 1254
rect -1410 1240 -1390 1254
rect -1390 1240 -1380 1254
rect -1360 1240 -1350 1254
rect -1350 1240 -1330 1254
rect -1330 1240 -1325 1254
rect -1305 1240 -1290 1254
rect -1290 1240 -1270 1254
rect -1470 1214 -1435 1220
rect -1415 1214 -1380 1220
rect -1360 1214 -1325 1220
rect -1305 1214 -1270 1220
rect -1470 1194 -1450 1214
rect -1450 1194 -1435 1214
rect -1415 1194 -1410 1214
rect -1410 1194 -1390 1214
rect -1390 1194 -1380 1214
rect -1360 1194 -1350 1214
rect -1350 1194 -1330 1214
rect -1330 1194 -1325 1214
rect -1305 1194 -1290 1214
rect -1290 1194 -1270 1214
rect -1470 1185 -1435 1194
rect -1415 1185 -1380 1194
rect -1360 1185 -1325 1194
rect -1305 1185 -1270 1194
rect -1085 1294 -1050 1305
rect -1030 1294 -995 1305
rect -975 1294 -940 1305
rect -920 1294 -885 1305
rect -1085 1274 -1070 1294
rect -1070 1274 -1050 1294
rect -1030 1274 -1010 1294
rect -1010 1274 -995 1294
rect -975 1274 -970 1294
rect -970 1274 -950 1294
rect -950 1274 -940 1294
rect -920 1274 -910 1294
rect -910 1274 -890 1294
rect -890 1274 -885 1294
rect -1085 1270 -1050 1274
rect -1030 1270 -995 1274
rect -975 1270 -940 1274
rect -920 1270 -885 1274
rect -1085 1234 -1070 1250
rect -1070 1234 -1050 1250
rect -1030 1234 -1010 1250
rect -1010 1234 -995 1250
rect -975 1234 -970 1250
rect -970 1234 -950 1250
rect -950 1234 -940 1250
rect -920 1234 -910 1250
rect -910 1234 -890 1250
rect -890 1234 -885 1250
rect -1085 1215 -1050 1234
rect -1030 1215 -995 1234
rect -975 1215 -940 1234
rect -920 1215 -885 1234
<< metal2 >>
rect -1095 1305 -875 1315
rect -1480 1275 -1260 1285
rect -1480 1240 -1470 1275
rect -1435 1240 -1415 1275
rect -1380 1240 -1360 1275
rect -1325 1240 -1305 1275
rect -1270 1240 -1260 1275
rect -1480 1220 -1260 1240
rect -1480 1185 -1470 1220
rect -1435 1185 -1415 1220
rect -1380 1185 -1360 1220
rect -1325 1185 -1305 1220
rect -1270 1185 -1260 1220
rect -1095 1270 -1085 1305
rect -1050 1270 -1030 1305
rect -995 1270 -975 1305
rect -940 1270 -920 1305
rect -885 1270 -875 1305
rect -1095 1250 -875 1270
rect -1095 1215 -1085 1250
rect -1050 1215 -1030 1250
rect -995 1215 -975 1250
rect -940 1215 -920 1250
rect -885 1215 -875 1250
rect -1095 1205 -875 1215
rect -1480 1175 -1260 1185
<< via2 >>
rect -1470 1240 -1435 1275
rect -1415 1240 -1380 1275
rect -1360 1240 -1325 1275
rect -1305 1240 -1270 1275
rect -1470 1185 -1435 1220
rect -1415 1185 -1380 1220
rect -1360 1185 -1325 1220
rect -1305 1185 -1270 1220
rect -1085 1270 -1050 1305
rect -1030 1270 -995 1305
rect -975 1270 -940 1305
rect -920 1270 -885 1305
rect -1085 1215 -1050 1250
rect -1030 1215 -995 1250
rect -975 1215 -940 1250
rect -920 1215 -885 1250
<< metal3 >>
rect -1095 1305 -875 1315
rect -1480 1275 -1260 1285
rect -1480 1240 -1470 1275
rect -1435 1240 -1415 1275
rect -1380 1240 -1360 1275
rect -1325 1240 -1305 1275
rect -1270 1240 -1260 1275
rect -1480 1220 -1260 1240
rect -1480 1185 -1470 1220
rect -1435 1185 -1415 1220
rect -1380 1185 -1360 1220
rect -1325 1185 -1305 1220
rect -1270 1185 -1260 1220
rect -1095 1270 -1085 1305
rect -1050 1270 -1030 1305
rect -995 1270 -975 1305
rect -940 1270 -920 1305
rect -885 1270 -875 1305
rect -1095 1250 -875 1270
rect -1095 1215 -1085 1250
rect -1050 1215 -1030 1250
rect -995 1215 -975 1250
rect -940 1215 -920 1250
rect -885 1215 -875 1250
rect -1095 1205 -875 1215
rect -1480 1175 -1260 1185
rect -1480 285 -675 1135
rect -1480 250 -1385 285
rect -1350 250 -1340 285
rect -1305 250 -1295 285
rect -1260 250 -1250 285
rect -1215 250 -1205 285
rect -1170 250 -1160 285
rect -1125 250 -1115 285
rect -1080 250 -1070 285
rect -1035 250 -1025 285
rect -990 250 -980 285
rect -945 250 -935 285
rect -900 250 -890 285
rect -855 250 -845 285
rect -810 250 -800 285
rect -765 250 -675 285
rect -1480 240 -675 250
rect -1480 205 -1385 240
rect -1350 205 -1340 240
rect -1305 205 -1295 240
rect -1260 205 -1250 240
rect -1215 205 -1205 240
rect -1170 205 -1160 240
rect -1125 205 -1115 240
rect -1080 205 -1070 240
rect -1035 205 -1025 240
rect -990 205 -980 240
rect -945 205 -935 240
rect -900 205 -890 240
rect -855 205 -845 240
rect -810 205 -800 240
rect -765 205 -675 240
rect -1480 195 -675 205
rect -1480 160 -1385 195
rect -1350 160 -1340 195
rect -1305 160 -1295 195
rect -1260 160 -1250 195
rect -1215 160 -1205 195
rect -1170 160 -1160 195
rect -1125 160 -1115 195
rect -1080 160 -1070 195
rect -1035 160 -1025 195
rect -990 160 -980 195
rect -945 160 -935 195
rect -900 160 -890 195
rect -855 160 -845 195
rect -810 160 -800 195
rect -765 160 -675 195
rect -1480 130 -675 160
<< via3 >>
rect -1470 1240 -1435 1275
rect -1415 1240 -1380 1275
rect -1360 1240 -1325 1275
rect -1305 1240 -1270 1275
rect -1470 1185 -1435 1220
rect -1415 1185 -1380 1220
rect -1360 1185 -1325 1220
rect -1305 1185 -1270 1220
rect -1085 1270 -1050 1305
rect -1030 1270 -995 1305
rect -975 1270 -940 1305
rect -920 1270 -885 1305
rect -1085 1215 -1050 1250
rect -1030 1215 -995 1250
rect -975 1215 -940 1250
rect -920 1215 -885 1250
rect -1385 250 -1350 285
rect -1340 250 -1305 285
rect -1295 250 -1260 285
rect -1250 250 -1215 285
rect -1205 250 -1170 285
rect -1160 250 -1125 285
rect -1115 250 -1080 285
rect -1070 250 -1035 285
rect -1025 250 -990 285
rect -980 250 -945 285
rect -935 250 -900 285
rect -890 250 -855 285
rect -845 250 -810 285
rect -800 250 -765 285
rect -1385 205 -1350 240
rect -1340 205 -1305 240
rect -1295 205 -1260 240
rect -1250 205 -1215 240
rect -1205 205 -1170 240
rect -1160 205 -1125 240
rect -1115 205 -1080 240
rect -1070 205 -1035 240
rect -1025 205 -990 240
rect -980 205 -945 240
rect -935 205 -900 240
rect -890 205 -855 240
rect -845 205 -810 240
rect -800 205 -765 240
rect -1385 160 -1350 195
rect -1340 160 -1305 195
rect -1295 160 -1260 195
rect -1250 160 -1215 195
rect -1205 160 -1170 195
rect -1160 160 -1125 195
rect -1115 160 -1080 195
rect -1070 160 -1035 195
rect -1025 160 -990 195
rect -980 160 -945 195
rect -935 160 -900 195
rect -890 160 -855 195
rect -845 160 -810 195
rect -800 160 -765 195
<< mimcap >>
rect -1465 1030 -690 1120
rect -1465 910 -1395 1030
rect -1275 910 -1230 1030
rect -1110 910 -1065 1030
rect -945 910 -900 1030
rect -780 910 -690 1030
rect -1465 865 -690 910
rect -1465 745 -1395 865
rect -1275 745 -1230 865
rect -1110 745 -1065 865
rect -945 745 -900 865
rect -780 745 -690 865
rect -1465 700 -690 745
rect -1465 580 -1395 700
rect -1275 580 -1230 700
rect -1110 580 -1065 700
rect -945 580 -900 700
rect -780 580 -690 700
rect -1465 535 -690 580
rect -1465 415 -1395 535
rect -1275 415 -1230 535
rect -1110 415 -1065 535
rect -945 415 -900 535
rect -780 415 -690 535
rect -1465 345 -690 415
<< mimcapcontact >>
rect -1395 910 -1275 1030
rect -1230 910 -1110 1030
rect -1065 910 -945 1030
rect -900 910 -780 1030
rect -1395 745 -1275 865
rect -1230 745 -1110 865
rect -1065 745 -945 865
rect -900 745 -780 865
rect -1395 580 -1275 700
rect -1230 580 -1110 700
rect -1065 580 -945 700
rect -900 580 -780 700
rect -1395 415 -1275 535
rect -1230 415 -1110 535
rect -1065 415 -945 535
rect -900 415 -780 535
<< metal4 >>
rect -1480 1275 -1240 1315
rect -1480 1240 -1470 1275
rect -1435 1240 -1415 1275
rect -1380 1240 -1360 1275
rect -1325 1240 -1305 1275
rect -1270 1240 -1240 1275
rect -1480 1220 -1240 1240
rect -1480 1185 -1470 1220
rect -1435 1185 -1415 1220
rect -1380 1185 -1360 1220
rect -1325 1185 -1305 1220
rect -1270 1185 -1240 1220
rect -1480 1135 -1240 1185
rect -1095 1305 -860 1350
rect -1095 1270 -1085 1305
rect -1050 1270 -1030 1305
rect -995 1270 -975 1305
rect -940 1270 -920 1305
rect -885 1270 -860 1305
rect -1095 1250 -860 1270
rect -1095 1215 -1085 1250
rect -1050 1215 -1030 1250
rect -995 1215 -975 1250
rect -940 1215 -920 1250
rect -885 1215 -860 1250
rect -1095 1175 -860 1215
rect -1480 1030 -675 1135
rect -1480 910 -1395 1030
rect -1275 910 -1230 1030
rect -1110 910 -1065 1030
rect -945 910 -900 1030
rect -780 910 -675 1030
rect -1480 865 -675 910
rect -1480 745 -1395 865
rect -1275 745 -1230 865
rect -1110 745 -1065 865
rect -945 745 -900 865
rect -780 745 -675 865
rect -1480 700 -675 745
rect -1480 580 -1395 700
rect -1275 580 -1230 700
rect -1110 580 -1065 700
rect -945 580 -900 700
rect -780 580 -675 700
rect -1480 535 -675 580
rect -1480 415 -1395 535
rect -1275 415 -1230 535
rect -1110 415 -1065 535
rect -945 415 -900 535
rect -780 415 -675 535
rect -1480 330 -675 415
rect -1405 285 -760 290
rect -1405 265 -1385 285
rect -1350 265 -1340 285
rect -1305 265 -1295 285
rect -1405 145 -1390 265
rect -1260 250 -1250 285
rect -1215 265 -1205 285
rect -1170 265 -1160 285
rect -1125 265 -1115 285
rect -1080 250 -1070 285
rect -1035 265 -1025 285
rect -990 265 -980 285
rect -945 265 -935 285
rect -940 250 -935 265
rect -900 265 -890 285
rect -855 265 -845 285
rect -810 265 -800 285
rect -900 250 -895 265
rect -765 250 -760 285
rect -1270 240 -1225 250
rect -1105 240 -1060 250
rect -940 240 -895 250
rect -775 240 -760 250
rect -1260 205 -1250 240
rect -1080 205 -1070 240
rect -940 205 -935 240
rect -900 205 -895 240
rect -765 205 -760 240
rect -1270 195 -1225 205
rect -1105 195 -1060 205
rect -940 195 -895 205
rect -775 195 -760 205
rect -1260 160 -1250 195
rect -1080 160 -1070 195
rect -940 160 -935 195
rect -900 160 -895 195
rect -765 160 -760 195
rect -1270 145 -1225 160
rect -1105 145 -1060 160
rect -940 145 -895 160
rect -775 145 -760 160
rect -1405 130 -760 145
<< via4 >>
rect -1390 250 -1385 265
rect -1385 250 -1350 265
rect -1350 250 -1340 265
rect -1340 250 -1305 265
rect -1305 250 -1295 265
rect -1295 250 -1270 265
rect -1225 250 -1215 265
rect -1215 250 -1205 265
rect -1205 250 -1170 265
rect -1170 250 -1160 265
rect -1160 250 -1125 265
rect -1125 250 -1115 265
rect -1115 250 -1105 265
rect -1060 250 -1035 265
rect -1035 250 -1025 265
rect -1025 250 -990 265
rect -990 250 -980 265
rect -980 250 -945 265
rect -945 250 -940 265
rect -895 250 -890 265
rect -890 250 -855 265
rect -855 250 -845 265
rect -845 250 -810 265
rect -810 250 -800 265
rect -800 250 -775 265
rect -1390 240 -1270 250
rect -1225 240 -1105 250
rect -1060 240 -940 250
rect -895 240 -775 250
rect -1390 205 -1385 240
rect -1385 205 -1350 240
rect -1350 205 -1340 240
rect -1340 205 -1305 240
rect -1305 205 -1295 240
rect -1295 205 -1270 240
rect -1225 205 -1215 240
rect -1215 205 -1205 240
rect -1205 205 -1170 240
rect -1170 205 -1160 240
rect -1160 205 -1125 240
rect -1125 205 -1115 240
rect -1115 205 -1105 240
rect -1060 205 -1035 240
rect -1035 205 -1025 240
rect -1025 205 -990 240
rect -990 205 -980 240
rect -980 205 -945 240
rect -945 205 -940 240
rect -895 205 -890 240
rect -890 205 -855 240
rect -855 205 -845 240
rect -845 205 -810 240
rect -810 205 -800 240
rect -800 205 -775 240
rect -1390 195 -1270 205
rect -1225 195 -1105 205
rect -1060 195 -940 205
rect -895 195 -775 205
rect -1390 160 -1385 195
rect -1385 160 -1350 195
rect -1350 160 -1340 195
rect -1340 160 -1305 195
rect -1305 160 -1295 195
rect -1295 160 -1270 195
rect -1225 160 -1215 195
rect -1215 160 -1205 195
rect -1205 160 -1170 195
rect -1170 160 -1160 195
rect -1160 160 -1125 195
rect -1125 160 -1115 195
rect -1115 160 -1105 195
rect -1060 160 -1035 195
rect -1035 160 -1025 195
rect -1025 160 -990 195
rect -990 160 -980 195
rect -980 160 -945 195
rect -945 160 -940 195
rect -895 160 -890 195
rect -890 160 -855 195
rect -855 160 -845 195
rect -845 160 -810 195
rect -810 160 -800 195
rect -800 160 -775 195
rect -1390 145 -1270 160
rect -1225 145 -1105 160
rect -1060 145 -940 160
rect -895 145 -775 160
<< mimcap2 >>
rect -1465 1030 -690 1120
rect -1465 910 -1395 1030
rect -1275 910 -1230 1030
rect -1110 910 -1065 1030
rect -945 910 -900 1030
rect -780 910 -690 1030
rect -1465 865 -690 910
rect -1465 745 -1395 865
rect -1275 745 -1230 865
rect -1110 745 -1065 865
rect -945 745 -900 865
rect -780 745 -690 865
rect -1465 700 -690 745
rect -1465 580 -1395 700
rect -1275 580 -1230 700
rect -1110 580 -1065 700
rect -945 580 -900 700
rect -780 580 -690 700
rect -1465 535 -690 580
rect -1465 415 -1395 535
rect -1275 415 -1230 535
rect -1110 415 -1065 535
rect -945 415 -900 535
rect -780 415 -690 535
rect -1465 345 -690 415
<< mimcap2contact >>
rect -1395 910 -1275 1030
rect -1230 910 -1110 1030
rect -1065 910 -945 1030
rect -900 910 -780 1030
rect -1395 745 -1275 865
rect -1230 745 -1110 865
rect -1065 745 -945 865
rect -900 745 -780 865
rect -1395 580 -1275 700
rect -1230 580 -1110 700
rect -1065 580 -945 700
rect -900 580 -780 700
rect -1395 415 -1275 535
rect -1230 415 -1110 535
rect -1065 415 -945 535
rect -900 415 -780 535
<< metal5 >>
rect -1480 1030 -675 1135
rect -1480 910 -1395 1030
rect -1275 910 -1230 1030
rect -1110 910 -1065 1030
rect -945 910 -900 1030
rect -780 910 -675 1030
rect -1480 865 -675 910
rect -1480 745 -1395 865
rect -1275 745 -1230 865
rect -1110 745 -1065 865
rect -945 745 -900 865
rect -780 745 -675 865
rect -1480 700 -675 745
rect -1480 580 -1395 700
rect -1275 580 -1230 700
rect -1110 580 -1065 700
rect -945 580 -900 700
rect -780 580 -675 700
rect -1480 535 -675 580
rect -1480 415 -1395 535
rect -1275 415 -1230 535
rect -1110 415 -1065 535
rect -945 415 -900 535
rect -780 415 -675 535
rect -1480 265 -675 415
rect -1480 145 -1390 265
rect -1270 145 -1225 265
rect -1105 145 -1060 265
rect -940 145 -895 265
rect -775 145 -675 265
rect -1480 130 -675 145
<< end >>
