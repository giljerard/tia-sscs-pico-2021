magic
tech sky130A
magscale 1 2
timestamp 1634930331
<< xpolycontact >>
rect -880 4130 -598 4610
rect -2220 -4898 -1938 -4420
rect -2220 -5660 -1938 -5180
rect 15380 4130 15662 4610
rect -330 -380 150 -98
rect 7150 -380 7630 -98
rect 14630 -380 15110 -98
rect -880 -6950 -598 -6470
rect 15380 -6950 15662 -6470
rect -2220 -8298 -1938 -7820
rect -2220 -9060 -1938 -8580
rect -270 -9900 210 -9618
rect 7210 -9900 7690 -9618
rect 14690 -9900 15170 -9618
<< xpolyres >>
rect -2220 -5180 -1938 -4898
rect -880 -6470 -598 4130
rect 150 -380 7150 -98
rect 7630 -380 14630 -98
rect 15380 -6470 15662 4130
rect -2220 -8580 -1938 -8298
rect 210 -9900 7210 -9618
rect 7690 -9900 14690 -9618
<< viali >>
rect -840 4550 -800 4590
rect -760 4550 -720 4590
rect -680 4550 -640 4590
rect -840 4470 -800 4510
rect -760 4470 -720 4510
rect -680 4470 -640 4510
rect -840 4390 -800 4430
rect -760 4390 -720 4430
rect -680 4390 -640 4430
rect -840 4310 -800 4350
rect -760 4310 -720 4350
rect -680 4310 -640 4350
rect -840 4230 -800 4270
rect -760 4230 -720 4270
rect -680 4230 -640 4270
rect -840 4150 -800 4190
rect -760 4150 -720 4190
rect -680 4150 -640 4190
rect 15420 4550 15460 4590
rect 15500 4550 15540 4590
rect 15580 4550 15620 4590
rect 15420 4470 15460 4510
rect 15500 4470 15540 4510
rect 15580 4470 15620 4510
rect 15420 4390 15460 4430
rect 15500 4390 15540 4430
rect 15580 4390 15620 4430
rect 15420 4310 15460 4350
rect 15500 4310 15540 4350
rect 15580 4310 15620 4350
rect 15420 4230 15460 4270
rect 15500 4230 15540 4270
rect 15580 4230 15620 4270
rect 15420 4150 15460 4190
rect 15500 4150 15540 4190
rect 15580 4150 15620 4190
rect -310 -180 -270 -140
rect -230 -180 -190 -140
rect -150 -180 -110 -140
rect -70 -180 -30 -140
rect 10 -180 50 -140
rect 90 -180 130 -140
rect -310 -260 -270 -220
rect -230 -260 -190 -220
rect -150 -260 -110 -220
rect -70 -260 -30 -220
rect 10 -260 50 -220
rect 90 -260 130 -220
rect -310 -340 -270 -300
rect -230 -340 -190 -300
rect -150 -340 -110 -300
rect -70 -340 -30 -300
rect 10 -340 50 -300
rect 90 -340 130 -300
rect 7170 -180 7210 -140
rect 7250 -180 7290 -140
rect 7330 -180 7370 -140
rect 7410 -180 7450 -140
rect 7490 -180 7530 -140
rect 7570 -180 7610 -140
rect 7170 -260 7210 -220
rect 7250 -260 7290 -220
rect 7330 -260 7370 -220
rect 7410 -260 7450 -220
rect 7490 -260 7530 -220
rect 7570 -260 7610 -220
rect 7170 -340 7210 -300
rect 7250 -340 7290 -300
rect 7330 -340 7370 -300
rect 7410 -340 7450 -300
rect 7490 -340 7530 -300
rect 7570 -340 7610 -300
rect 14650 -180 14690 -140
rect 14730 -180 14770 -140
rect 14810 -180 14850 -140
rect 14890 -180 14930 -140
rect 14970 -180 15010 -140
rect 15050 -180 15090 -140
rect 14650 -260 14690 -220
rect 14730 -260 14770 -220
rect 14810 -260 14850 -220
rect 14890 -260 14930 -220
rect 14970 -260 15010 -220
rect 15050 -260 15090 -220
rect 14650 -340 14690 -300
rect 14730 -340 14770 -300
rect 14810 -340 14850 -300
rect 14890 -340 14930 -300
rect 14970 -340 15010 -300
rect 15050 -340 15090 -300
rect -2178 -4480 -2138 -4440
rect -2098 -4480 -2058 -4440
rect -2018 -4480 -1978 -4440
rect -2178 -4560 -2138 -4520
rect -2098 -4560 -2058 -4520
rect -2018 -4560 -1978 -4520
rect -2178 -4640 -2138 -4600
rect -2098 -4640 -2058 -4600
rect -2018 -4640 -1978 -4600
rect -2178 -4720 -2138 -4680
rect -2098 -4720 -2058 -4680
rect -2018 -4720 -1978 -4680
rect -2178 -4800 -2138 -4760
rect -2098 -4800 -2058 -4760
rect -2018 -4800 -1978 -4760
rect -2178 -4880 -2138 -4840
rect -2098 -4880 -2058 -4840
rect -2018 -4880 -1978 -4840
rect -2178 -5240 -2138 -5200
rect -2098 -5240 -2058 -5200
rect -2018 -5240 -1978 -5200
rect -2178 -5320 -2138 -5280
rect -2098 -5320 -2058 -5280
rect -2018 -5320 -1978 -5280
rect -2178 -5400 -2138 -5360
rect -2098 -5400 -2058 -5360
rect -2018 -5400 -1978 -5360
rect -2178 -5480 -2138 -5440
rect -2098 -5480 -2058 -5440
rect -2018 -5480 -1978 -5440
rect -2178 -5560 -2138 -5520
rect -2098 -5560 -2058 -5520
rect -2018 -5560 -1978 -5520
rect -2178 -5640 -2138 -5600
rect -2098 -5640 -2058 -5600
rect -2018 -5640 -1978 -5600
rect -840 -6530 -800 -6490
rect -760 -6530 -720 -6490
rect -680 -6530 -640 -6490
rect -840 -6610 -800 -6570
rect -760 -6610 -720 -6570
rect -680 -6610 -640 -6570
rect -840 -6690 -800 -6650
rect -760 -6690 -720 -6650
rect -680 -6690 -640 -6650
rect -840 -6770 -800 -6730
rect -760 -6770 -720 -6730
rect -680 -6770 -640 -6730
rect -840 -6850 -800 -6810
rect -760 -6850 -720 -6810
rect -680 -6850 -640 -6810
rect -840 -6930 -800 -6890
rect -760 -6930 -720 -6890
rect -680 -6930 -640 -6890
rect 15420 -6530 15460 -6490
rect 15500 -6530 15540 -6490
rect 15580 -6530 15620 -6490
rect 15420 -6610 15460 -6570
rect 15500 -6610 15540 -6570
rect 15580 -6610 15620 -6570
rect 15420 -6690 15460 -6650
rect 15500 -6690 15540 -6650
rect 15580 -6690 15620 -6650
rect 15420 -6770 15460 -6730
rect 15500 -6770 15540 -6730
rect 15580 -6770 15620 -6730
rect 15420 -6850 15460 -6810
rect 15500 -6850 15540 -6810
rect 15580 -6850 15620 -6810
rect 15420 -6930 15460 -6890
rect 15500 -6930 15540 -6890
rect 15580 -6930 15620 -6890
rect -2178 -7880 -2138 -7840
rect -2098 -7880 -2058 -7840
rect -2018 -7880 -1978 -7840
rect -2178 -7960 -2138 -7920
rect -2098 -7960 -2058 -7920
rect -2018 -7960 -1978 -7920
rect -2178 -8040 -2138 -8000
rect -2098 -8040 -2058 -8000
rect -2018 -8040 -1978 -8000
rect -2178 -8120 -2138 -8080
rect -2098 -8120 -2058 -8080
rect -2018 -8120 -1978 -8080
rect -2178 -8200 -2138 -8160
rect -2098 -8200 -2058 -8160
rect -2018 -8200 -1978 -8160
rect -2178 -8280 -2138 -8240
rect -2098 -8280 -2058 -8240
rect -2018 -8280 -1978 -8240
rect -2178 -8640 -2138 -8600
rect -2098 -8640 -2058 -8600
rect -2018 -8640 -1978 -8600
rect -2178 -8720 -2138 -8680
rect -2098 -8720 -2058 -8680
rect -2018 -8720 -1978 -8680
rect -2178 -8800 -2138 -8760
rect -2098 -8800 -2058 -8760
rect -2018 -8800 -1978 -8760
rect -2178 -8880 -2138 -8840
rect -2098 -8880 -2058 -8840
rect -2018 -8880 -1978 -8840
rect -2178 -8960 -2138 -8920
rect -2098 -8960 -2058 -8920
rect -2018 -8960 -1978 -8920
rect -2178 -9040 -2138 -9000
rect -2098 -9040 -2058 -9000
rect -2018 -9040 -1978 -9000
rect -250 -9700 -210 -9660
rect -170 -9700 -130 -9660
rect -90 -9700 -50 -9660
rect -10 -9700 30 -9660
rect 70 -9700 110 -9660
rect 150 -9700 190 -9660
rect -250 -9780 -210 -9740
rect -170 -9780 -130 -9740
rect -90 -9780 -50 -9740
rect -10 -9780 30 -9740
rect 70 -9780 110 -9740
rect 150 -9780 190 -9740
rect -250 -9860 -210 -9820
rect -170 -9860 -130 -9820
rect -90 -9860 -50 -9820
rect -10 -9860 30 -9820
rect 70 -9860 110 -9820
rect 150 -9860 190 -9820
rect 7230 -9700 7270 -9660
rect 7310 -9700 7350 -9660
rect 7390 -9700 7430 -9660
rect 7470 -9700 7510 -9660
rect 7550 -9700 7590 -9660
rect 7630 -9700 7670 -9660
rect 7230 -9780 7270 -9740
rect 7310 -9780 7350 -9740
rect 7390 -9780 7430 -9740
rect 7470 -9780 7510 -9740
rect 7550 -9780 7590 -9740
rect 7630 -9780 7670 -9740
rect 7230 -9860 7270 -9820
rect 7310 -9860 7350 -9820
rect 7390 -9860 7430 -9820
rect 7470 -9860 7510 -9820
rect 7550 -9860 7590 -9820
rect 7630 -9860 7670 -9820
rect 14710 -9700 14750 -9660
rect 14790 -9700 14830 -9660
rect 14870 -9700 14910 -9660
rect 14950 -9700 14990 -9660
rect 15030 -9700 15070 -9660
rect 15110 -9700 15150 -9660
rect 14710 -9780 14750 -9740
rect 14790 -9780 14830 -9740
rect 14870 -9780 14910 -9740
rect 14950 -9780 14990 -9740
rect 15030 -9780 15070 -9740
rect 15110 -9780 15150 -9740
rect 14710 -9860 14750 -9820
rect 14790 -9860 14830 -9820
rect 14870 -9860 14910 -9820
rect 14950 -9860 14990 -9820
rect 15030 -9860 15070 -9820
rect 15110 -9860 15150 -9820
<< metal1 >>
rect 21060 7210 21540 7230
rect 21060 7140 21090 7210
rect 21160 7140 21200 7210
rect 21270 7140 21310 7210
rect 21380 7140 21420 7210
rect 21490 7140 21540 7210
rect 21060 7100 21540 7140
rect 21060 7030 21090 7100
rect 21160 7030 21200 7100
rect 21270 7030 21310 7100
rect 21380 7030 21420 7100
rect 21490 7030 21540 7100
rect 21060 6920 21540 7030
rect 23460 7210 23940 7230
rect 23460 7140 23490 7210
rect 23560 7140 23600 7210
rect 23670 7140 23710 7210
rect 23780 7140 23820 7210
rect 23890 7140 23940 7210
rect 23460 7100 23940 7140
rect 23460 7030 23490 7100
rect 23560 7030 23600 7100
rect 23670 7030 23710 7100
rect 23780 7030 23820 7100
rect 23890 7030 23940 7100
rect 23460 6950 23940 7030
rect 11760 6880 13360 6900
rect 1540 6850 3140 6870
rect 1540 6780 1570 6850
rect 1640 6780 1680 6850
rect 1750 6780 1790 6850
rect 1860 6780 1900 6850
rect 1970 6780 2010 6850
rect 2080 6780 2120 6850
rect 2190 6780 2230 6850
rect 2300 6780 2340 6850
rect 2410 6780 2450 6850
rect 2520 6780 2560 6850
rect 2630 6780 2670 6850
rect 2740 6780 2780 6850
rect 2850 6780 2890 6850
rect 2960 6780 3000 6850
rect 3070 6780 3140 6850
rect 1540 6740 3140 6780
rect 1540 6670 1570 6740
rect 1640 6670 1680 6740
rect 1750 6670 1790 6740
rect 1860 6670 1900 6740
rect 1970 6670 2010 6740
rect 2080 6670 2120 6740
rect 2190 6670 2230 6740
rect 2300 6670 2340 6740
rect 2410 6670 2450 6740
rect 2520 6670 2560 6740
rect 2630 6670 2670 6740
rect 2740 6670 2780 6740
rect 2850 6670 2890 6740
rect 2960 6670 3000 6740
rect 3070 6670 3140 6740
rect 1540 6520 3140 6670
rect 11760 6810 11790 6880
rect 11860 6810 11900 6880
rect 11970 6810 12010 6880
rect 12080 6810 12120 6880
rect 12190 6810 12230 6880
rect 12300 6810 12340 6880
rect 12410 6810 12450 6880
rect 12520 6810 12560 6880
rect 12630 6810 12670 6880
rect 12740 6810 12780 6880
rect 12850 6810 12890 6880
rect 12960 6810 13000 6880
rect 13070 6810 13110 6880
rect 13180 6810 13220 6880
rect 13290 6810 13360 6880
rect 11760 6770 13360 6810
rect 11760 6700 11790 6770
rect 11860 6700 11900 6770
rect 11970 6700 12010 6770
rect 12080 6700 12120 6770
rect 12190 6700 12230 6770
rect 12300 6700 12340 6770
rect 12410 6700 12450 6770
rect 12520 6700 12560 6770
rect 12630 6700 12670 6770
rect 12740 6700 12780 6770
rect 12850 6700 12890 6770
rect 12960 6700 13000 6770
rect 13070 6700 13110 6770
rect 13180 6700 13220 6770
rect 13290 6700 13360 6770
rect 11760 6550 13360 6700
rect 7400 5390 7490 5410
rect 7400 5320 7410 5390
rect 7480 5320 7490 5390
rect 7400 5280 7490 5320
rect 7400 5210 7410 5280
rect 7480 5210 7490 5280
rect 7400 5170 7490 5210
rect 7400 5100 7410 5170
rect 7480 5100 7490 5170
rect 7400 5060 7490 5100
rect 7400 4990 7410 5060
rect 7480 4990 7490 5060
rect 7400 4950 7490 4990
rect 7400 4880 7410 4950
rect 7480 4880 7490 4950
rect 7400 4860 7490 4880
rect -880 4590 -598 4610
rect -880 4390 -840 4590
rect -800 4580 -760 4590
rect -770 4550 -760 4580
rect -720 4580 -680 4590
rect -720 4550 -710 4580
rect -770 4510 -710 4550
rect -800 4470 -760 4510
rect -720 4470 -680 4510
rect -770 4430 -710 4470
rect -770 4400 -760 4430
rect -800 4390 -760 4400
rect -720 4400 -710 4430
rect -720 4390 -680 4400
rect -640 4390 -598 4590
rect -880 4360 -598 4390
rect -880 4290 -840 4360
rect -770 4350 -710 4360
rect -770 4310 -760 4350
rect -720 4310 -710 4350
rect -770 4290 -710 4310
rect -640 4290 -598 4360
rect -880 4270 -598 4290
rect -880 4150 -840 4270
rect -800 4250 -760 4270
rect -770 4230 -760 4250
rect -720 4250 -680 4270
rect -720 4230 -710 4250
rect -770 4190 -710 4230
rect -770 4180 -760 4190
rect -800 4150 -760 4180
rect -720 4180 -710 4190
rect -720 4150 -680 4180
rect -640 4150 -598 4270
rect -880 4130 -598 4150
rect 15380 4590 15662 4610
rect 15380 4390 15420 4590
rect 15460 4580 15500 4590
rect 15490 4550 15500 4580
rect 15540 4580 15580 4590
rect 15540 4550 15550 4580
rect 15490 4510 15550 4550
rect 15460 4470 15500 4510
rect 15540 4470 15580 4510
rect 15490 4430 15550 4470
rect 15490 4400 15500 4430
rect 15460 4390 15500 4400
rect 15540 4400 15550 4430
rect 15540 4390 15580 4400
rect 15620 4390 15662 4590
rect 15380 4360 15662 4390
rect 15380 4290 15420 4360
rect 15490 4350 15550 4360
rect 15490 4310 15500 4350
rect 15540 4310 15550 4350
rect 15490 4290 15550 4310
rect 15620 4290 15662 4360
rect 15380 4270 15662 4290
rect 15380 4150 15420 4270
rect 15460 4250 15500 4270
rect 15490 4230 15500 4250
rect 15540 4250 15580 4270
rect 15540 4230 15550 4250
rect 15490 4190 15550 4230
rect 15490 4180 15500 4190
rect 15460 4150 15500 4180
rect 15540 4180 15550 4190
rect 15540 4150 15580 4180
rect 15620 4150 15662 4270
rect 15380 4130 15662 4150
rect 19400 3990 19720 5440
rect 22300 3360 22630 3380
rect 22300 3290 22320 3360
rect 22390 3290 22430 3360
rect 22500 3290 22540 3360
rect 22610 3290 22630 3360
rect 22300 3250 22630 3290
rect 22300 3180 22320 3250
rect 22390 3180 22430 3250
rect 22500 3180 22540 3250
rect 22610 3180 22630 3250
rect 22300 3140 22630 3180
rect 22300 3070 22320 3140
rect 22390 3070 22430 3140
rect 22500 3070 22540 3140
rect 22610 3070 22630 3140
rect 22300 3050 22630 3070
rect 20020 2600 20500 2670
rect 20020 2530 20070 2600
rect 20140 2530 20180 2600
rect 20250 2530 20290 2600
rect 20360 2530 20400 2600
rect 20470 2530 20500 2600
rect 20020 2490 20500 2530
rect 20020 2420 20070 2490
rect 20140 2420 20180 2490
rect 20250 2420 20290 2490
rect 20360 2420 20400 2490
rect 20470 2420 20500 2490
rect 20020 2400 20500 2420
rect 24500 2600 24980 2660
rect 24500 2530 24550 2600
rect 24620 2530 24660 2600
rect 24730 2530 24770 2600
rect 24840 2530 24880 2600
rect 24950 2530 24980 2600
rect 24500 2490 24980 2530
rect 24500 2420 24550 2490
rect 24620 2420 24660 2490
rect 24730 2420 24770 2490
rect 24840 2420 24880 2490
rect 24950 2420 24980 2490
rect 24500 2400 24980 2420
rect 14590 1160 14900 1180
rect 14590 1090 14600 1160
rect 14670 1090 14700 1160
rect 14770 1090 14810 1160
rect 14880 1090 14900 1160
rect 14590 1050 14900 1090
rect 14590 980 14600 1050
rect 14670 980 14700 1050
rect 14770 980 14810 1050
rect 14880 980 14900 1050
rect 14590 940 14900 980
rect 14590 870 14600 940
rect 14670 870 14700 940
rect 14770 870 14810 940
rect 14880 870 14900 940
rect 14590 850 14900 870
rect 21060 920 21540 940
rect 21060 850 21090 920
rect 21160 850 21200 920
rect 21270 850 21310 920
rect 21380 850 21420 920
rect 21490 850 21540 920
rect 21060 810 21540 850
rect 21060 740 21090 810
rect 21160 740 21200 810
rect 21270 740 21310 810
rect 21380 740 21420 810
rect 21490 740 21540 810
rect 21060 640 21540 740
rect 23460 920 23940 940
rect 23460 850 23490 920
rect 23560 850 23600 920
rect 23670 850 23710 920
rect 23780 850 23820 920
rect 23890 850 23940 920
rect 23460 810 23940 850
rect 23460 740 23490 810
rect 23560 740 23600 810
rect 23670 740 23710 810
rect 23780 740 23820 810
rect 23890 740 23940 810
rect 23460 650 23940 740
rect -330 -140 150 -98
rect -330 -180 -310 -140
rect -110 -180 -80 -140
rect -10 -180 10 -140
rect 130 -180 150 -140
rect -330 -210 -300 -180
rect -230 -210 -190 -180
rect -120 -210 -80 -180
rect -10 -210 30 -180
rect 100 -210 150 -180
rect -330 -220 150 -210
rect -330 -260 -310 -220
rect -270 -260 -230 -220
rect -190 -260 -150 -220
rect -110 -260 -70 -220
rect -30 -260 10 -220
rect 50 -260 90 -220
rect 130 -260 150 -220
rect -330 -270 150 -260
rect -330 -300 -300 -270
rect -230 -300 -190 -270
rect -120 -300 -80 -270
rect -10 -300 30 -270
rect 100 -300 150 -270
rect -330 -340 -310 -300
rect -110 -340 -80 -300
rect -10 -340 10 -300
rect 130 -340 150 -300
rect -330 -380 150 -340
rect 1080 -790 2680 40
rect 7150 -120 7630 -98
rect 7150 -140 7180 -120
rect 7240 -140 7280 -120
rect 7340 -140 7440 -120
rect 7500 -140 7540 -120
rect 7600 -140 7630 -120
rect 7150 -180 7170 -140
rect 7240 -180 7250 -140
rect 7370 -180 7410 -140
rect 7530 -180 7540 -140
rect 7610 -180 7630 -140
rect 7150 -210 7630 -180
rect 7150 -220 7180 -210
rect 7240 -220 7280 -210
rect 7340 -220 7440 -210
rect 7500 -220 7540 -210
rect 7600 -220 7630 -210
rect 7150 -260 7170 -220
rect 7240 -260 7250 -220
rect 7370 -260 7410 -220
rect 7530 -260 7540 -220
rect 7610 -260 7630 -220
rect 7150 -270 7180 -260
rect 7240 -270 7280 -260
rect 7340 -270 7440 -260
rect 7500 -270 7540 -260
rect 7600 -270 7630 -260
rect 7150 -300 7630 -270
rect 7150 -340 7170 -300
rect 7240 -340 7250 -300
rect 7370 -340 7410 -300
rect 7530 -340 7540 -300
rect 7610 -340 7630 -300
rect 7150 -360 7180 -340
rect 7240 -360 7280 -340
rect 7340 -360 7440 -340
rect 7500 -360 7540 -340
rect 7600 -360 7630 -340
rect 7150 -380 7630 -360
rect 1080 -860 1150 -790
rect 1220 -860 1260 -790
rect 1330 -860 1370 -790
rect 1440 -860 1480 -790
rect 1550 -860 1590 -790
rect 1660 -860 1700 -790
rect 1770 -860 1810 -790
rect 1880 -860 1920 -790
rect 1990 -860 2030 -790
rect 2100 -860 2140 -790
rect 2210 -860 2250 -790
rect 2320 -860 2360 -790
rect 2430 -860 2470 -790
rect 2540 -860 2580 -790
rect 2650 -860 2680 -790
rect 1080 -900 2680 -860
rect 1080 -970 1150 -900
rect 1220 -970 1260 -900
rect 1330 -970 1370 -900
rect 1440 -970 1480 -900
rect 1550 -970 1590 -900
rect 1660 -970 1700 -900
rect 1770 -970 1810 -900
rect 1880 -970 1920 -900
rect 1990 -970 2030 -900
rect 2100 -970 2140 -900
rect 2210 -970 2250 -900
rect 2320 -970 2360 -900
rect 2430 -970 2470 -900
rect 2540 -970 2580 -900
rect 2650 -970 2680 -900
rect 1080 -990 2680 -970
rect 12220 -790 13820 40
rect 14630 -140 15110 -98
rect 14630 -180 14650 -140
rect 14850 -180 14880 -140
rect 14950 -180 14970 -140
rect 15090 -180 15110 -140
rect 14630 -210 14660 -180
rect 14730 -210 14770 -180
rect 14840 -210 14880 -180
rect 14950 -210 14990 -180
rect 15060 -210 15110 -180
rect 14630 -220 15110 -210
rect 14630 -260 14650 -220
rect 14690 -260 14730 -220
rect 14770 -260 14810 -220
rect 14850 -260 14890 -220
rect 14930 -260 14970 -220
rect 15010 -260 15050 -220
rect 15090 -260 15110 -220
rect 14630 -270 15110 -260
rect 14630 -300 14660 -270
rect 14730 -300 14770 -270
rect 14840 -300 14880 -270
rect 14950 -300 14990 -270
rect 15060 -300 15110 -270
rect 14630 -340 14650 -300
rect 14850 -340 14880 -300
rect 14950 -340 14970 -300
rect 15090 -340 15110 -300
rect 14630 -380 15110 -340
rect 12220 -860 12250 -790
rect 12320 -860 12360 -790
rect 12430 -860 12470 -790
rect 12540 -860 12580 -790
rect 12650 -860 12690 -790
rect 12760 -860 12800 -790
rect 12870 -860 12910 -790
rect 12980 -860 13020 -790
rect 13090 -860 13130 -790
rect 13200 -860 13240 -790
rect 13310 -860 13350 -790
rect 13420 -860 13460 -790
rect 13530 -860 13570 -790
rect 13640 -860 13680 -790
rect 13750 -860 13820 -790
rect 12220 -900 13820 -860
rect 12220 -970 12250 -900
rect 12320 -970 12360 -900
rect 12430 -970 12470 -900
rect 12540 -970 12580 -900
rect 12650 -970 12690 -900
rect 12760 -970 12800 -900
rect 12870 -970 12910 -900
rect 12980 -970 13020 -900
rect 13090 -970 13130 -900
rect 13200 -970 13240 -900
rect 13310 -970 13350 -900
rect 13420 -970 13460 -900
rect 13530 -970 13570 -900
rect 13640 -970 13680 -900
rect 13750 -970 13820 -900
rect 12220 -990 13820 -970
rect 19400 -2040 19660 -820
rect 1540 -2780 3140 -2760
rect 1540 -2850 1570 -2780
rect 1640 -2850 1680 -2780
rect 1750 -2850 1790 -2780
rect 1860 -2850 1900 -2780
rect 1970 -2850 2010 -2780
rect 2080 -2850 2120 -2780
rect 2190 -2850 2230 -2780
rect 2300 -2850 2340 -2780
rect 2410 -2850 2450 -2780
rect 2520 -2850 2560 -2780
rect 2630 -2850 2670 -2780
rect 2740 -2850 2780 -2780
rect 2850 -2850 2890 -2780
rect 2960 -2850 3000 -2780
rect 3070 -2850 3140 -2780
rect 1540 -2890 3140 -2850
rect 1540 -2960 1570 -2890
rect 1640 -2960 1680 -2890
rect 1750 -2960 1790 -2890
rect 1860 -2960 1900 -2890
rect 1970 -2960 2010 -2890
rect 2080 -2960 2120 -2890
rect 2190 -2960 2230 -2890
rect 2300 -2960 2340 -2890
rect 2410 -2960 2450 -2890
rect 2520 -2960 2560 -2890
rect 2630 -2960 2670 -2890
rect 2740 -2960 2780 -2890
rect 2850 -2960 2890 -2890
rect 2960 -2960 3000 -2890
rect 3070 -2960 3140 -2890
rect 1540 -3020 3140 -2960
rect 11760 -2780 13360 -2760
rect 11760 -2850 11790 -2780
rect 11860 -2850 11900 -2780
rect 11970 -2850 12010 -2780
rect 12080 -2850 12120 -2780
rect 12190 -2850 12230 -2780
rect 12300 -2850 12340 -2780
rect 12410 -2850 12450 -2780
rect 12520 -2850 12560 -2780
rect 12630 -2850 12670 -2780
rect 12740 -2850 12780 -2780
rect 12850 -2850 12890 -2780
rect 12960 -2850 13000 -2780
rect 13070 -2850 13110 -2780
rect 13180 -2850 13220 -2780
rect 13290 -2850 13360 -2780
rect 11760 -2890 13360 -2850
rect 11760 -2960 11790 -2890
rect 11860 -2960 11900 -2890
rect 11970 -2960 12010 -2890
rect 12080 -2960 12120 -2890
rect 12190 -2960 12230 -2890
rect 12300 -2960 12340 -2890
rect 12410 -2960 12450 -2890
rect 12520 -2960 12560 -2890
rect 12630 -2960 12670 -2890
rect 12740 -2960 12780 -2890
rect 12850 -2960 12890 -2890
rect 12960 -2960 13000 -2890
rect 13070 -2960 13110 -2890
rect 13180 -2960 13220 -2890
rect 13290 -2960 13360 -2890
rect 11760 -3020 13360 -2960
rect 22320 -3050 22650 -3030
rect 22320 -3120 22340 -3050
rect 22410 -3120 22450 -3050
rect 22520 -3120 22560 -3050
rect 22630 -3120 22650 -3050
rect 22320 -3160 22650 -3120
rect 22320 -3230 22340 -3160
rect 22410 -3230 22450 -3160
rect 22520 -3230 22560 -3160
rect 22630 -3230 22650 -3160
rect 22320 -3270 22650 -3230
rect 22320 -3340 22340 -3270
rect 22410 -3340 22450 -3270
rect 22520 -3340 22560 -3270
rect 22630 -3340 22650 -3270
rect 22320 -3360 22650 -3340
rect 20020 -3690 20500 -3630
rect 20020 -3760 20070 -3690
rect 20140 -3760 20180 -3690
rect 20250 -3760 20290 -3690
rect 20360 -3760 20400 -3690
rect 20470 -3760 20500 -3690
rect 20020 -3800 20500 -3760
rect 20020 -3870 20070 -3800
rect 20140 -3870 20180 -3800
rect 20250 -3870 20290 -3800
rect 20360 -3870 20400 -3800
rect 20470 -3870 20500 -3800
rect 20020 -3890 20500 -3870
rect 24500 -3690 24980 -3630
rect 24500 -3760 24550 -3690
rect 24620 -3760 24660 -3690
rect 24730 -3760 24770 -3690
rect 24840 -3760 24880 -3690
rect 24950 -3760 24980 -3690
rect 24500 -3800 24980 -3760
rect 24500 -3870 24550 -3800
rect 24620 -3870 24660 -3800
rect 24730 -3870 24770 -3800
rect 24840 -3870 24880 -3800
rect 24950 -3870 24980 -3800
rect 24500 -3890 24980 -3870
rect -2220 -4440 -1938 -4420
rect -2220 -4470 -2178 -4440
rect -2138 -4470 -2098 -4440
rect -2058 -4470 -2018 -4440
rect -2220 -4540 -2200 -4470
rect -2130 -4480 -2098 -4470
rect -2020 -4480 -2018 -4470
rect -1978 -4480 -1938 -4440
rect -2130 -4520 -2090 -4480
rect -2020 -4520 -1938 -4480
rect -2130 -4540 -2098 -4520
rect -2020 -4540 -2018 -4520
rect -2220 -4560 -2178 -4540
rect -2138 -4560 -2098 -4540
rect -2058 -4560 -2018 -4540
rect -1978 -4560 -1938 -4520
rect -2220 -4580 -1938 -4560
rect -2220 -4650 -2200 -4580
rect -2130 -4600 -2090 -4580
rect -2020 -4600 -1938 -4580
rect -2130 -4640 -2098 -4600
rect -2020 -4640 -2018 -4600
rect -1978 -4640 -1938 -4600
rect -2130 -4650 -2090 -4640
rect -2020 -4650 -1938 -4640
rect -2220 -4680 -1938 -4650
rect -2220 -4690 -2178 -4680
rect -2138 -4690 -2098 -4680
rect -2058 -4690 -2018 -4680
rect -2220 -4760 -2200 -4690
rect -2130 -4720 -2098 -4690
rect -2020 -4720 -2018 -4690
rect -1978 -4720 -1938 -4680
rect -2130 -4760 -2090 -4720
rect -2020 -4760 -1938 -4720
rect -2220 -4800 -2178 -4760
rect -2138 -4800 -2098 -4760
rect -2058 -4800 -2018 -4760
rect -1978 -4800 -1938 -4760
rect -2220 -4870 -2200 -4800
rect -2130 -4840 -2090 -4800
rect -2020 -4840 -1938 -4800
rect -2130 -4870 -2098 -4840
rect -2020 -4870 -2018 -4840
rect -2220 -4880 -2178 -4870
rect -2138 -4880 -2098 -4870
rect -2058 -4880 -2018 -4870
rect -1978 -4880 -1938 -4840
rect 7290 -4560 7620 -4540
rect 7290 -4630 7310 -4560
rect 7380 -4630 7420 -4560
rect 7490 -4630 7530 -4560
rect 7600 -4630 7620 -4560
rect 7290 -4670 7620 -4630
rect 7290 -4740 7310 -4670
rect 7380 -4740 7420 -4670
rect 7490 -4740 7530 -4670
rect 7600 -4740 7620 -4670
rect 7290 -4780 7620 -4740
rect 7290 -4850 7310 -4780
rect 7380 -4850 7420 -4780
rect 7490 -4850 7530 -4780
rect 7600 -4850 7620 -4780
rect 7290 -4870 7620 -4850
rect -2220 -4898 -1938 -4880
rect -2220 -5200 -1938 -5180
rect -2220 -5240 -2178 -5200
rect -2138 -5240 -2098 -5200
rect -2058 -5240 -2018 -5200
rect -1978 -5240 -1938 -5200
rect -2220 -5280 -2140 -5240
rect -2070 -5280 -2030 -5240
rect -2220 -5320 -2178 -5280
rect -2058 -5310 -2030 -5280
rect -1960 -5310 -1938 -5240
rect -2138 -5320 -2098 -5310
rect -2058 -5320 -2018 -5310
rect -1978 -5320 -1938 -5310
rect -2220 -5350 -1938 -5320
rect -2220 -5360 -2140 -5350
rect -2070 -5360 -2030 -5350
rect -2220 -5400 -2178 -5360
rect -2058 -5400 -2030 -5360
rect -2220 -5420 -2140 -5400
rect -2070 -5420 -2030 -5400
rect -1960 -5420 -1938 -5350
rect -2220 -5440 -1938 -5420
rect -2220 -5480 -2178 -5440
rect -2138 -5460 -2098 -5440
rect -2058 -5460 -2018 -5440
rect -1978 -5460 -1938 -5440
rect -2058 -5480 -2030 -5460
rect -2220 -5520 -2140 -5480
rect -2070 -5520 -2030 -5480
rect -2220 -5560 -2178 -5520
rect -2058 -5530 -2030 -5520
rect -1960 -5530 -1938 -5460
rect -2138 -5560 -2098 -5530
rect -2058 -5560 -2018 -5530
rect -1978 -5560 -1938 -5530
rect -2220 -5570 -1938 -5560
rect -2220 -5600 -2140 -5570
rect -2070 -5600 -2030 -5570
rect -2220 -5640 -2178 -5600
rect -2058 -5640 -2030 -5600
rect -1960 -5640 -1938 -5570
rect -2220 -5660 -1938 -5640
rect 7570 -6460 7870 -6420
rect -880 -6490 -598 -6470
rect -880 -6690 -840 -6490
rect -800 -6500 -760 -6490
rect -770 -6530 -760 -6500
rect -720 -6500 -680 -6490
rect -720 -6530 -710 -6500
rect -770 -6570 -710 -6530
rect -800 -6610 -760 -6570
rect -720 -6610 -680 -6570
rect -770 -6650 -710 -6610
rect -770 -6680 -760 -6650
rect -800 -6690 -760 -6680
rect -720 -6680 -710 -6650
rect -720 -6690 -680 -6680
rect -640 -6690 -598 -6490
rect 7570 -6520 7590 -6460
rect 7650 -6520 7690 -6460
rect 7750 -6520 7790 -6460
rect 7850 -6520 7870 -6460
rect 7570 -6560 7870 -6520
rect 7570 -6620 7590 -6560
rect 7650 -6620 7690 -6560
rect 7750 -6620 7790 -6560
rect 7850 -6620 7870 -6560
rect 7570 -6660 7870 -6620
rect -880 -6720 -598 -6690
rect -880 -6790 -840 -6720
rect -770 -6730 -710 -6720
rect -770 -6770 -760 -6730
rect -720 -6770 -710 -6730
rect -770 -6790 -710 -6770
rect -640 -6790 -598 -6720
rect 7570 -6720 7590 -6660
rect 7650 -6720 7690 -6660
rect 7750 -6720 7790 -6660
rect 7850 -6720 7870 -6660
rect 15380 -6490 15662 -6470
rect 7570 -6760 7870 -6720
rect 15380 -6690 15420 -6490
rect 15460 -6500 15500 -6490
rect 15490 -6530 15500 -6500
rect 15540 -6500 15580 -6490
rect 15540 -6530 15550 -6500
rect 15490 -6570 15550 -6530
rect 15460 -6610 15500 -6570
rect 15540 -6610 15580 -6570
rect 15490 -6650 15550 -6610
rect 15490 -6680 15500 -6650
rect 15460 -6690 15500 -6680
rect 15540 -6680 15550 -6650
rect 15540 -6690 15580 -6680
rect 15620 -6690 15662 -6490
rect 15380 -6720 15662 -6690
rect -880 -6810 -598 -6790
rect -880 -6930 -840 -6810
rect -800 -6830 -760 -6810
rect -770 -6850 -760 -6830
rect -720 -6830 -680 -6810
rect -720 -6850 -710 -6830
rect -770 -6890 -710 -6850
rect -770 -6900 -760 -6890
rect -800 -6930 -760 -6900
rect -720 -6900 -710 -6890
rect -720 -6930 -680 -6900
rect -640 -6930 -598 -6810
rect 7570 -6820 7590 -6760
rect 7650 -6820 7690 -6760
rect 7750 -6820 7790 -6760
rect 7850 -6820 7870 -6760
rect 7570 -6850 7870 -6820
rect 15380 -6790 15420 -6720
rect 15490 -6730 15550 -6720
rect 15490 -6770 15500 -6730
rect 15540 -6770 15550 -6730
rect 15490 -6790 15550 -6770
rect 15620 -6790 15662 -6720
rect 15380 -6810 15662 -6790
rect 15380 -6930 15420 -6810
rect 15460 -6830 15500 -6810
rect 15490 -6850 15500 -6830
rect 15540 -6830 15580 -6810
rect 15540 -6850 15550 -6830
rect 15490 -6890 15550 -6850
rect 15490 -6900 15500 -6890
rect 15460 -6930 15500 -6900
rect 15540 -6900 15550 -6890
rect 15540 -6930 15580 -6900
rect 15620 -6930 15662 -6810
rect -880 -6950 -598 -6930
rect 15380 -6950 15662 -6930
rect -2220 -7840 -1938 -7820
rect -2220 -7870 -2178 -7840
rect -2138 -7870 -2098 -7840
rect -2058 -7870 -2018 -7840
rect -2220 -7940 -2200 -7870
rect -2130 -7880 -2098 -7870
rect -2020 -7880 -2018 -7870
rect -1978 -7880 -1938 -7840
rect -2130 -7920 -2090 -7880
rect -2020 -7920 -1938 -7880
rect -2130 -7940 -2098 -7920
rect -2020 -7940 -2018 -7920
rect -2220 -7960 -2178 -7940
rect -2138 -7960 -2098 -7940
rect -2058 -7960 -2018 -7940
rect -1978 -7960 -1938 -7920
rect -2220 -7980 -1938 -7960
rect -2220 -8050 -2200 -7980
rect -2130 -8000 -2090 -7980
rect -2020 -8000 -1938 -7980
rect -2130 -8040 -2098 -8000
rect -2020 -8040 -2018 -8000
rect -1978 -8040 -1938 -8000
rect -2130 -8050 -2090 -8040
rect -2020 -8050 -1938 -8040
rect -2220 -8080 -1938 -8050
rect -2220 -8090 -2178 -8080
rect -2138 -8090 -2098 -8080
rect -2058 -8090 -2018 -8080
rect -2220 -8160 -2200 -8090
rect -2130 -8120 -2098 -8090
rect -2020 -8120 -2018 -8090
rect -1978 -8120 -1938 -8080
rect -2130 -8160 -2090 -8120
rect -2020 -8160 -1938 -8120
rect -2220 -8200 -2178 -8160
rect -2138 -8200 -2098 -8160
rect -2058 -8200 -2018 -8160
rect -1978 -8200 -1938 -8160
rect -2220 -8270 -2200 -8200
rect -2130 -8240 -2090 -8200
rect -2020 -8240 -1938 -8200
rect -2130 -8270 -2098 -8240
rect -2020 -8270 -2018 -8240
rect -2220 -8280 -2178 -8270
rect -2138 -8280 -2098 -8270
rect -2058 -8280 -2018 -8270
rect -1978 -8280 -1938 -8240
rect -2220 -8298 -1938 -8280
rect 14590 -8230 14900 -8210
rect 14590 -8300 14600 -8230
rect 14670 -8300 14700 -8230
rect 14770 -8300 14810 -8230
rect 14880 -8300 14900 -8230
rect 14590 -8340 14900 -8300
rect 14590 -8410 14600 -8340
rect 14670 -8410 14700 -8340
rect 14770 -8410 14810 -8340
rect 14880 -8410 14900 -8340
rect 14590 -8450 14900 -8410
rect 14590 -8520 14600 -8450
rect 14670 -8520 14700 -8450
rect 14770 -8520 14810 -8450
rect 14880 -8520 14900 -8450
rect 14590 -8540 14900 -8520
rect 19210 -8560 20140 -8530
rect -2220 -8600 -1938 -8580
rect -2220 -8640 -2178 -8600
rect -2138 -8640 -2098 -8600
rect -2058 -8640 -2018 -8600
rect -1978 -8640 -1938 -8600
rect -2220 -8680 -2140 -8640
rect -2070 -8680 -2030 -8640
rect -2220 -8720 -2178 -8680
rect -2058 -8710 -2030 -8680
rect -1960 -8710 -1938 -8640
rect -2138 -8720 -2098 -8710
rect -2058 -8720 -2018 -8710
rect -1978 -8720 -1938 -8710
rect -2220 -8750 -1938 -8720
rect -2220 -8760 -2140 -8750
rect -2070 -8760 -2030 -8750
rect -2220 -8800 -2178 -8760
rect -2058 -8800 -2030 -8760
rect -2220 -8820 -2140 -8800
rect -2070 -8820 -2030 -8800
rect -1960 -8820 -1938 -8750
rect -2220 -8840 -1938 -8820
rect -2220 -8880 -2178 -8840
rect -2138 -8860 -2098 -8840
rect -2058 -8860 -2018 -8840
rect -1978 -8860 -1938 -8840
rect 19210 -8630 19230 -8560
rect 19300 -8630 19330 -8560
rect 19400 -8630 19430 -8560
rect 19500 -8630 20140 -8560
rect 19210 -8660 20140 -8630
rect 19210 -8730 19230 -8660
rect 19300 -8730 19330 -8660
rect 19400 -8730 19430 -8660
rect 19500 -8730 20140 -8660
rect 19210 -8760 20140 -8730
rect 19210 -8830 19230 -8760
rect 19300 -8830 19330 -8760
rect 19400 -8830 19430 -8760
rect 19500 -8830 20140 -8760
rect 19210 -8850 20140 -8830
rect -2058 -8880 -2030 -8860
rect -2220 -8920 -2140 -8880
rect -2070 -8920 -2030 -8880
rect -2220 -8960 -2178 -8920
rect -2058 -8930 -2030 -8920
rect -1960 -8930 -1938 -8860
rect -2138 -8960 -2098 -8930
rect -2058 -8960 -2018 -8930
rect -1978 -8960 -1938 -8930
rect -2220 -8970 -1938 -8960
rect -2220 -9000 -2140 -8970
rect -2070 -9000 -2030 -8970
rect -2220 -9040 -2178 -9000
rect -2058 -9040 -2030 -9000
rect -1960 -9040 -1938 -8970
rect -2220 -9060 -1938 -9040
rect 19940 -9000 20260 -8970
rect 19940 -9070 19960 -9000
rect 20030 -9070 20060 -9000
rect 20130 -9070 20160 -9000
rect 20230 -9070 20260 -9000
rect 19940 -9100 20260 -9070
rect 19940 -9170 19960 -9100
rect 20030 -9170 20060 -9100
rect 20130 -9170 20160 -9100
rect 20230 -9170 20260 -9100
rect 19940 -9200 20260 -9170
rect 19940 -9270 19960 -9200
rect 20030 -9270 20060 -9200
rect 20130 -9270 20160 -9200
rect 20230 -9270 20260 -9200
rect 19940 -9290 20260 -9270
rect -270 -9660 210 -9618
rect -270 -9700 -250 -9660
rect -50 -9700 -20 -9660
rect 50 -9700 70 -9660
rect 190 -9700 210 -9660
rect -270 -9730 -240 -9700
rect -170 -9730 -130 -9700
rect -60 -9730 -20 -9700
rect 50 -9730 90 -9700
rect 160 -9730 210 -9700
rect -270 -9740 210 -9730
rect -270 -9780 -250 -9740
rect -210 -9780 -170 -9740
rect -130 -9780 -90 -9740
rect -50 -9780 -10 -9740
rect 30 -9780 70 -9740
rect 110 -9780 150 -9740
rect 190 -9780 210 -9740
rect -270 -9790 210 -9780
rect -270 -9820 -240 -9790
rect -170 -9820 -130 -9790
rect -60 -9820 -20 -9790
rect 50 -9820 90 -9790
rect 160 -9820 210 -9790
rect -270 -9860 -250 -9820
rect -50 -9860 -20 -9820
rect 50 -9860 70 -9820
rect 190 -9860 210 -9820
rect -270 -9900 210 -9860
rect 1080 -10340 2680 -9500
rect 7210 -9640 7690 -9618
rect 7210 -9660 7240 -9640
rect 7300 -9660 7340 -9640
rect 7400 -9660 7500 -9640
rect 7560 -9660 7600 -9640
rect 7660 -9660 7690 -9640
rect 7210 -9700 7230 -9660
rect 7300 -9700 7310 -9660
rect 7430 -9700 7470 -9660
rect 7590 -9700 7600 -9660
rect 7670 -9700 7690 -9660
rect 7210 -9730 7690 -9700
rect 7210 -9740 7240 -9730
rect 7300 -9740 7340 -9730
rect 7400 -9740 7500 -9730
rect 7560 -9740 7600 -9730
rect 7660 -9740 7690 -9730
rect 7210 -9780 7230 -9740
rect 7300 -9780 7310 -9740
rect 7430 -9780 7470 -9740
rect 7590 -9780 7600 -9740
rect 7670 -9780 7690 -9740
rect 7210 -9790 7240 -9780
rect 7300 -9790 7340 -9780
rect 7400 -9790 7500 -9780
rect 7560 -9790 7600 -9780
rect 7660 -9790 7690 -9780
rect 7210 -9820 7690 -9790
rect 7210 -9860 7230 -9820
rect 7300 -9860 7310 -9820
rect 7430 -9860 7470 -9820
rect 7590 -9860 7600 -9820
rect 7670 -9860 7690 -9820
rect 7210 -9880 7240 -9860
rect 7300 -9880 7340 -9860
rect 7400 -9880 7500 -9860
rect 7560 -9880 7600 -9860
rect 7660 -9880 7690 -9860
rect 7210 -9900 7690 -9880
rect 1080 -10410 1150 -10340
rect 1220 -10410 1260 -10340
rect 1330 -10410 1370 -10340
rect 1440 -10410 1480 -10340
rect 1550 -10410 1590 -10340
rect 1660 -10410 1700 -10340
rect 1770 -10410 1810 -10340
rect 1880 -10410 1920 -10340
rect 1990 -10410 2030 -10340
rect 2100 -10410 2140 -10340
rect 2210 -10410 2250 -10340
rect 2320 -10410 2360 -10340
rect 2430 -10410 2470 -10340
rect 2540 -10410 2580 -10340
rect 2650 -10410 2680 -10340
rect 1080 -10450 2680 -10410
rect 1080 -10520 1150 -10450
rect 1220 -10520 1260 -10450
rect 1330 -10520 1370 -10450
rect 1440 -10520 1480 -10450
rect 1550 -10520 1590 -10450
rect 1660 -10520 1700 -10450
rect 1770 -10520 1810 -10450
rect 1880 -10520 1920 -10450
rect 1990 -10520 2030 -10450
rect 2100 -10520 2140 -10450
rect 2210 -10520 2250 -10450
rect 2320 -10520 2360 -10450
rect 2430 -10520 2470 -10450
rect 2540 -10520 2580 -10450
rect 2650 -10520 2680 -10450
rect 1080 -10540 2680 -10520
rect 12220 -10370 13820 -9520
rect 14690 -9660 15170 -9618
rect 14690 -9700 14710 -9660
rect 14910 -9700 14940 -9660
rect 15010 -9700 15030 -9660
rect 15150 -9700 15170 -9660
rect 14690 -9730 14720 -9700
rect 14790 -9730 14830 -9700
rect 14900 -9730 14940 -9700
rect 15010 -9730 15050 -9700
rect 15120 -9730 15170 -9700
rect 14690 -9740 15170 -9730
rect 14690 -9780 14710 -9740
rect 14750 -9780 14790 -9740
rect 14830 -9780 14870 -9740
rect 14910 -9780 14950 -9740
rect 14990 -9780 15030 -9740
rect 15070 -9780 15110 -9740
rect 15150 -9780 15170 -9740
rect 14690 -9790 15170 -9780
rect 14690 -9820 14720 -9790
rect 14790 -9820 14830 -9790
rect 14900 -9820 14940 -9790
rect 15010 -9820 15050 -9790
rect 15120 -9820 15170 -9790
rect 14690 -9860 14710 -9820
rect 14910 -9860 14940 -9820
rect 15010 -9860 15030 -9820
rect 15150 -9860 15170 -9820
rect 14690 -9900 15170 -9860
rect 12220 -10440 12290 -10370
rect 12360 -10440 12400 -10370
rect 12470 -10440 12510 -10370
rect 12580 -10440 12620 -10370
rect 12690 -10440 12730 -10370
rect 12800 -10440 12840 -10370
rect 12910 -10440 12950 -10370
rect 13020 -10440 13060 -10370
rect 13130 -10440 13170 -10370
rect 13240 -10440 13280 -10370
rect 13350 -10440 13390 -10370
rect 13460 -10440 13500 -10370
rect 13570 -10440 13610 -10370
rect 13680 -10440 13720 -10370
rect 13790 -10440 13820 -10370
rect 12220 -10480 13820 -10440
rect 12220 -10550 12290 -10480
rect 12360 -10550 12400 -10480
rect 12470 -10550 12510 -10480
rect 12580 -10550 12620 -10480
rect 12690 -10550 12730 -10480
rect 12800 -10550 12840 -10480
rect 12910 -10550 12950 -10480
rect 13020 -10550 13060 -10480
rect 13130 -10550 13170 -10480
rect 13240 -10550 13280 -10480
rect 13350 -10550 13390 -10480
rect 13460 -10550 13500 -10480
rect 13570 -10550 13610 -10480
rect 13680 -10550 13720 -10480
rect 13790 -10550 13820 -10480
rect 12220 -10570 13820 -10550
rect 2210 -12300 3810 -12280
rect 2210 -12370 2240 -12300
rect 2310 -12370 2350 -12300
rect 2420 -12370 2460 -12300
rect 2530 -12370 2570 -12300
rect 2640 -12370 2680 -12300
rect 2750 -12370 2790 -12300
rect 2860 -12370 2900 -12300
rect 2970 -12370 3010 -12300
rect 3080 -12370 3120 -12300
rect 3190 -12370 3230 -12300
rect 3300 -12370 3340 -12300
rect 3410 -12370 3450 -12300
rect 3520 -12370 3560 -12300
rect 3630 -12370 3670 -12300
rect 3740 -12370 3810 -12300
rect 2210 -12410 3810 -12370
rect 2210 -12480 2240 -12410
rect 2310 -12480 2350 -12410
rect 2420 -12480 2460 -12410
rect 2530 -12480 2570 -12410
rect 2640 -12480 2680 -12410
rect 2750 -12480 2790 -12410
rect 2860 -12480 2900 -12410
rect 2970 -12480 3010 -12410
rect 3080 -12480 3120 -12410
rect 3190 -12480 3230 -12410
rect 3300 -12480 3340 -12410
rect 3410 -12480 3450 -12410
rect 3520 -12480 3560 -12410
rect 3630 -12480 3670 -12410
rect 3740 -12480 3810 -12410
rect 2210 -12550 3810 -12480
rect 11090 -12300 12690 -12280
rect 11090 -12370 11120 -12300
rect 11190 -12370 11230 -12300
rect 11300 -12370 11340 -12300
rect 11410 -12370 11450 -12300
rect 11520 -12370 11560 -12300
rect 11630 -12370 11670 -12300
rect 11740 -12370 11780 -12300
rect 11850 -12370 11890 -12300
rect 11960 -12370 12000 -12300
rect 12070 -12370 12110 -12300
rect 12180 -12370 12220 -12300
rect 12290 -12370 12330 -12300
rect 12400 -12370 12440 -12300
rect 12510 -12370 12550 -12300
rect 12620 -12370 12690 -12300
rect 11090 -12410 12690 -12370
rect 11090 -12480 11120 -12410
rect 11190 -12480 11230 -12410
rect 11300 -12480 11340 -12410
rect 11410 -12480 11450 -12410
rect 11520 -12480 11560 -12410
rect 11630 -12480 11670 -12410
rect 11740 -12480 11780 -12410
rect 11850 -12480 11890 -12410
rect 11960 -12480 12000 -12410
rect 12070 -12480 12110 -12410
rect 12180 -12480 12220 -12410
rect 12290 -12480 12330 -12410
rect 12400 -12480 12440 -12410
rect 12510 -12480 12550 -12410
rect 12620 -12480 12690 -12410
rect 11090 -12550 12690 -12480
rect 19210 -14220 20420 -14190
rect 19210 -14290 19230 -14220
rect 19300 -14290 19330 -14220
rect 19400 -14290 19430 -14220
rect 19500 -14290 20420 -14220
rect 19210 -14320 20420 -14290
rect 19210 -14390 19230 -14320
rect 19300 -14390 19330 -14320
rect 19400 -14390 19430 -14320
rect 19500 -14390 20420 -14320
rect 19210 -14420 20420 -14390
rect 19210 -14490 19230 -14420
rect 19300 -14490 19330 -14420
rect 19400 -14490 19430 -14420
rect 19500 -14490 20420 -14420
rect 19210 -14510 20420 -14490
rect 20460 -14870 20780 -14840
rect 20460 -14940 20480 -14870
rect 20550 -14940 20580 -14870
rect 20650 -14940 20680 -14870
rect 20750 -14940 20780 -14870
rect 20460 -14970 20780 -14940
rect 20460 -15040 20480 -14970
rect 20550 -15040 20580 -14970
rect 20650 -15040 20680 -14970
rect 20750 -15040 20780 -14970
rect 20460 -15070 20780 -15040
rect 20460 -15140 20480 -15070
rect 20550 -15140 20580 -15070
rect 20650 -15140 20680 -15070
rect 20750 -15140 20780 -15070
rect 20460 -15160 20780 -15140
rect 7210 -17600 7650 -17580
rect 7210 -17670 7230 -17600
rect 7300 -17670 7340 -17600
rect 7410 -17670 7450 -17600
rect 7520 -17670 7560 -17600
rect 7630 -17670 7650 -17600
rect 7210 -17710 7650 -17670
rect 7210 -17780 7230 -17710
rect 7300 -17780 7340 -17710
rect 7410 -17780 7450 -17710
rect 7520 -17780 7560 -17710
rect 7630 -17780 7650 -17710
rect 7210 -17820 7650 -17780
rect 7210 -17890 7230 -17820
rect 7300 -17890 7340 -17820
rect 7410 -17890 7450 -17820
rect 7520 -17890 7560 -17820
rect 7630 -17890 7650 -17820
rect 7210 -17930 7650 -17890
rect 7210 -18000 7230 -17930
rect 7300 -18000 7340 -17930
rect 7410 -18000 7450 -17930
rect 7520 -18000 7560 -17930
rect 7630 -18000 7650 -17930
rect 7210 -18020 7650 -18000
rect 19210 -20290 20220 -20260
rect 19210 -20360 19230 -20290
rect 19300 -20360 19330 -20290
rect 19400 -20360 19430 -20290
rect 19500 -20360 20220 -20290
rect 19210 -20390 20220 -20360
rect 19210 -20460 19230 -20390
rect 19300 -20460 19330 -20390
rect 19400 -20460 19430 -20390
rect 19500 -20460 20220 -20390
rect 19210 -20490 20220 -20460
rect 19210 -20560 19230 -20490
rect 19300 -20560 19330 -20490
rect 19400 -20560 19430 -20490
rect 19500 -20560 20220 -20490
rect 19210 -20580 20220 -20560
rect 20020 -20720 20340 -20690
rect 20020 -20790 20040 -20720
rect 20110 -20790 20140 -20720
rect 20210 -20790 20240 -20720
rect 20310 -20790 20340 -20720
rect 20020 -20820 20340 -20790
rect 20020 -20890 20040 -20820
rect 20110 -20890 20140 -20820
rect 20210 -20890 20240 -20820
rect 20310 -20890 20340 -20820
rect 20020 -20920 20340 -20890
rect 20020 -20990 20040 -20920
rect 20110 -20990 20140 -20920
rect 20210 -20990 20240 -20920
rect 20310 -20990 20340 -20920
rect 20020 -21010 20340 -20990
rect 2210 -22660 3810 -22590
rect 2210 -22730 2280 -22660
rect 2350 -22730 2390 -22660
rect 2460 -22730 2500 -22660
rect 2570 -22730 2610 -22660
rect 2680 -22730 2720 -22660
rect 2790 -22730 2830 -22660
rect 2900 -22730 2940 -22660
rect 3010 -22730 3050 -22660
rect 3120 -22730 3160 -22660
rect 3230 -22730 3270 -22660
rect 3340 -22730 3380 -22660
rect 3450 -22730 3490 -22660
rect 3560 -22730 3600 -22660
rect 3670 -22730 3710 -22660
rect 3780 -22730 3810 -22660
rect 2210 -22770 3810 -22730
rect 2210 -22840 2280 -22770
rect 2350 -22840 2390 -22770
rect 2460 -22840 2500 -22770
rect 2570 -22840 2610 -22770
rect 2680 -22840 2720 -22770
rect 2790 -22840 2830 -22770
rect 2900 -22840 2940 -22770
rect 3010 -22840 3050 -22770
rect 3120 -22840 3160 -22770
rect 3230 -22840 3270 -22770
rect 3340 -22840 3380 -22770
rect 3450 -22840 3490 -22770
rect 3560 -22840 3600 -22770
rect 3670 -22840 3710 -22770
rect 3780 -22840 3810 -22770
rect 2210 -22860 3810 -22840
rect 11090 -22660 12690 -22590
rect 11090 -22730 11160 -22660
rect 11230 -22730 11270 -22660
rect 11340 -22730 11380 -22660
rect 11450 -22730 11490 -22660
rect 11560 -22730 11600 -22660
rect 11670 -22730 11710 -22660
rect 11780 -22730 11820 -22660
rect 11890 -22730 11930 -22660
rect 12000 -22730 12040 -22660
rect 12110 -22730 12150 -22660
rect 12220 -22730 12260 -22660
rect 12330 -22730 12370 -22660
rect 12440 -22730 12480 -22660
rect 12550 -22730 12590 -22660
rect 12660 -22730 12690 -22660
rect 11090 -22770 12690 -22730
rect 11090 -22840 11160 -22770
rect 11230 -22840 11270 -22770
rect 11340 -22840 11380 -22770
rect 11450 -22840 11490 -22770
rect 11560 -22840 11600 -22770
rect 11670 -22840 11710 -22770
rect 11780 -22840 11820 -22770
rect 11890 -22840 11930 -22770
rect 12000 -22840 12040 -22770
rect 12110 -22840 12150 -22770
rect 12220 -22840 12260 -22770
rect 12330 -22840 12370 -22770
rect 12440 -22840 12480 -22770
rect 12550 -22840 12590 -22770
rect 12660 -22840 12690 -22770
rect 11090 -22860 12690 -22840
<< via1 >>
rect 21090 7140 21160 7210
rect 21200 7140 21270 7210
rect 21310 7140 21380 7210
rect 21420 7140 21490 7210
rect 21090 7030 21160 7100
rect 21200 7030 21270 7100
rect 21310 7030 21380 7100
rect 21420 7030 21490 7100
rect 23490 7140 23560 7210
rect 23600 7140 23670 7210
rect 23710 7140 23780 7210
rect 23820 7140 23890 7210
rect 23490 7030 23560 7100
rect 23600 7030 23670 7100
rect 23710 7030 23780 7100
rect 23820 7030 23890 7100
rect 1570 6780 1640 6850
rect 1680 6780 1750 6850
rect 1790 6780 1860 6850
rect 1900 6780 1970 6850
rect 2010 6780 2080 6850
rect 2120 6780 2190 6850
rect 2230 6780 2300 6850
rect 2340 6780 2410 6850
rect 2450 6780 2520 6850
rect 2560 6780 2630 6850
rect 2670 6780 2740 6850
rect 2780 6780 2850 6850
rect 2890 6780 2960 6850
rect 3000 6780 3070 6850
rect 1570 6670 1640 6740
rect 1680 6670 1750 6740
rect 1790 6670 1860 6740
rect 1900 6670 1970 6740
rect 2010 6670 2080 6740
rect 2120 6670 2190 6740
rect 2230 6670 2300 6740
rect 2340 6670 2410 6740
rect 2450 6670 2520 6740
rect 2560 6670 2630 6740
rect 2670 6670 2740 6740
rect 2780 6670 2850 6740
rect 2890 6670 2960 6740
rect 3000 6670 3070 6740
rect 11790 6810 11860 6880
rect 11900 6810 11970 6880
rect 12010 6810 12080 6880
rect 12120 6810 12190 6880
rect 12230 6810 12300 6880
rect 12340 6810 12410 6880
rect 12450 6810 12520 6880
rect 12560 6810 12630 6880
rect 12670 6810 12740 6880
rect 12780 6810 12850 6880
rect 12890 6810 12960 6880
rect 13000 6810 13070 6880
rect 13110 6810 13180 6880
rect 13220 6810 13290 6880
rect 11790 6700 11860 6770
rect 11900 6700 11970 6770
rect 12010 6700 12080 6770
rect 12120 6700 12190 6770
rect 12230 6700 12300 6770
rect 12340 6700 12410 6770
rect 12450 6700 12520 6770
rect 12560 6700 12630 6770
rect 12670 6700 12740 6770
rect 12780 6700 12850 6770
rect 12890 6700 12960 6770
rect 13000 6700 13070 6770
rect 13110 6700 13180 6770
rect 13220 6700 13290 6770
rect 7380 6230 7440 6290
rect 7480 6230 7540 6290
rect 20380 6210 20450 6280
rect 20490 6210 20560 6280
rect 20600 6210 20670 6280
rect 20710 6210 20780 6280
rect 7380 6080 7440 6190
rect 7480 6080 7540 6190
rect 20380 6100 20450 6170
rect 20490 6100 20560 6170
rect 20600 6100 20670 6170
rect 20710 6100 20780 6170
rect 7380 5980 7440 6040
rect 7480 5980 7540 6040
rect 20380 5990 20450 6060
rect 20490 5990 20560 6060
rect 20600 5990 20670 6060
rect 20710 5990 20780 6060
rect 7410 5320 7480 5390
rect 7410 5210 7480 5280
rect 7410 5100 7480 5170
rect 7410 4990 7480 5060
rect 7410 4880 7480 4950
rect -840 4550 -800 4580
rect -800 4550 -770 4580
rect -710 4550 -680 4580
rect -680 4550 -640 4580
rect -840 4510 -770 4550
rect -710 4510 -640 4550
rect -840 4430 -770 4470
rect -710 4430 -640 4470
rect -840 4400 -800 4430
rect -800 4400 -770 4430
rect -710 4400 -680 4430
rect -680 4400 -640 4430
rect -840 4350 -770 4360
rect -710 4350 -640 4360
rect -840 4310 -800 4350
rect -800 4310 -770 4350
rect -710 4310 -680 4350
rect -680 4310 -640 4350
rect -840 4290 -770 4310
rect -710 4290 -640 4310
rect -840 4230 -800 4250
rect -800 4230 -770 4250
rect -710 4230 -680 4250
rect -680 4230 -640 4250
rect -840 4190 -770 4230
rect -710 4190 -640 4230
rect -840 4180 -800 4190
rect -800 4180 -770 4190
rect -710 4180 -680 4190
rect -680 4180 -640 4190
rect 15420 4550 15460 4580
rect 15460 4550 15490 4580
rect 15550 4550 15580 4580
rect 15580 4550 15620 4580
rect 15420 4510 15490 4550
rect 15550 4510 15620 4550
rect 15420 4430 15490 4470
rect 15550 4430 15620 4470
rect 15420 4400 15460 4430
rect 15460 4400 15490 4430
rect 15550 4400 15580 4430
rect 15580 4400 15620 4430
rect 15420 4350 15490 4360
rect 15550 4350 15620 4360
rect 15420 4310 15460 4350
rect 15460 4310 15490 4350
rect 15550 4310 15580 4350
rect 15580 4310 15620 4350
rect 15420 4290 15490 4310
rect 15550 4290 15620 4310
rect 15420 4230 15460 4250
rect 15460 4230 15490 4250
rect 15550 4230 15580 4250
rect 15580 4230 15620 4250
rect 15420 4190 15490 4230
rect 15550 4190 15620 4230
rect 15420 4180 15460 4190
rect 15460 4180 15490 4190
rect 15550 4180 15580 4190
rect 15580 4180 15620 4190
rect 25310 4810 25370 4870
rect 25410 4810 25470 4870
rect 25510 4810 25570 4870
rect 25310 4710 25370 4770
rect 25410 4710 25470 4770
rect 25510 4710 25570 4770
rect 25310 4610 25370 4670
rect 25410 4610 25470 4670
rect 25510 4610 25570 4670
rect 25310 4510 25370 4570
rect 25410 4510 25470 4570
rect 25510 4510 25570 4570
rect 25310 4410 25370 4470
rect 25410 4410 25470 4470
rect 25510 4410 25570 4470
rect 25310 4310 25370 4370
rect 25410 4310 25470 4370
rect 25510 4310 25570 4370
rect 25310 4210 25370 4270
rect 25410 4210 25470 4270
rect 25510 4210 25570 4270
rect 25310 4110 25370 4170
rect 25410 4110 25470 4170
rect 25510 4110 25570 4170
rect 25310 4010 25370 4070
rect 25410 4010 25470 4070
rect 25510 4010 25570 4070
rect 22320 3290 22390 3360
rect 22430 3290 22500 3360
rect 22540 3290 22610 3360
rect 7050 3180 7110 3240
rect 7150 3180 7210 3240
rect 7250 3180 7310 3240
rect 7590 3180 7650 3240
rect 7690 3180 7750 3240
rect 7790 3180 7850 3240
rect 22320 3180 22390 3250
rect 22430 3180 22500 3250
rect 22540 3180 22610 3250
rect 7050 3080 7110 3140
rect 7150 3080 7210 3140
rect 7250 3080 7310 3140
rect 7590 3080 7650 3140
rect 7690 3080 7750 3140
rect 7790 3080 7850 3140
rect 22320 3070 22390 3140
rect 22430 3070 22500 3140
rect 22540 3070 22610 3140
rect 7050 2980 7110 3040
rect 7150 2980 7210 3040
rect 7250 2980 7310 3040
rect 7590 2980 7650 3040
rect 7690 2980 7750 3040
rect 7790 2980 7850 3040
rect 4770 2830 4830 2890
rect 4870 2830 4930 2890
rect 4970 2830 5030 2890
rect 9870 2830 9930 2890
rect 9970 2830 10030 2890
rect 10070 2830 10130 2890
rect 4770 2730 4830 2790
rect 4870 2730 4930 2790
rect 4970 2730 5030 2790
rect 9870 2730 9930 2790
rect 9970 2730 10030 2790
rect 10070 2730 10130 2790
rect 4770 2630 4830 2690
rect 4870 2630 4930 2690
rect 4970 2630 5030 2690
rect 9870 2630 9930 2690
rect 9970 2630 10030 2690
rect 10070 2630 10130 2690
rect 20070 2530 20140 2600
rect 20180 2530 20250 2600
rect 20290 2530 20360 2600
rect 20400 2530 20470 2600
rect 20070 2420 20140 2490
rect 20180 2420 20250 2490
rect 20290 2420 20360 2490
rect 20400 2420 20470 2490
rect 24550 2530 24620 2600
rect 24660 2530 24730 2600
rect 24770 2530 24840 2600
rect 24880 2530 24950 2600
rect 24550 2420 24620 2490
rect 24660 2420 24730 2490
rect 24770 2420 24840 2490
rect 24880 2420 24950 2490
rect 14600 1090 14670 1160
rect 14700 1090 14770 1160
rect 14810 1090 14880 1160
rect 14600 980 14670 1050
rect 14700 980 14770 1050
rect 14810 980 14880 1050
rect 14600 870 14670 940
rect 14700 870 14770 940
rect 14810 870 14880 940
rect 21090 850 21160 920
rect 21200 850 21270 920
rect 21310 850 21380 920
rect 21420 850 21490 920
rect 21090 740 21160 810
rect 21200 740 21270 810
rect 21310 740 21380 810
rect 21420 740 21490 810
rect 23490 850 23560 920
rect 23600 850 23670 920
rect 23710 850 23780 920
rect 23820 850 23890 920
rect 23490 740 23560 810
rect 23600 740 23670 810
rect 23710 740 23780 810
rect 23820 740 23890 810
rect -300 -180 -270 -140
rect -270 -180 -230 -140
rect -190 -180 -150 -140
rect -150 -180 -120 -140
rect -80 -180 -70 -140
rect -70 -180 -30 -140
rect -30 -180 -10 -140
rect 30 -180 50 -140
rect 50 -180 90 -140
rect 90 -180 100 -140
rect -300 -210 -230 -180
rect -190 -210 -120 -180
rect -80 -210 -10 -180
rect 30 -210 100 -180
rect -300 -300 -230 -270
rect -190 -300 -120 -270
rect -80 -300 -10 -270
rect 30 -300 100 -270
rect -300 -340 -270 -300
rect -270 -340 -230 -300
rect -190 -340 -150 -300
rect -150 -340 -120 -300
rect -80 -340 -70 -300
rect -70 -340 -30 -300
rect -30 -340 -10 -300
rect 30 -340 50 -300
rect 50 -340 90 -300
rect 90 -340 100 -300
rect 7180 -140 7240 -120
rect 7280 -140 7340 -120
rect 7440 -140 7500 -120
rect 7540 -140 7600 -120
rect 7180 -180 7210 -140
rect 7210 -180 7240 -140
rect 7280 -180 7290 -140
rect 7290 -180 7330 -140
rect 7330 -180 7340 -140
rect 7440 -180 7450 -140
rect 7450 -180 7490 -140
rect 7490 -180 7500 -140
rect 7540 -180 7570 -140
rect 7570 -180 7600 -140
rect 7180 -220 7240 -210
rect 7280 -220 7340 -210
rect 7440 -220 7500 -210
rect 7540 -220 7600 -210
rect 7180 -260 7210 -220
rect 7210 -260 7240 -220
rect 7280 -260 7290 -220
rect 7290 -260 7330 -220
rect 7330 -260 7340 -220
rect 7440 -260 7450 -220
rect 7450 -260 7490 -220
rect 7490 -260 7500 -220
rect 7540 -260 7570 -220
rect 7570 -260 7600 -220
rect 7180 -270 7240 -260
rect 7280 -270 7340 -260
rect 7440 -270 7500 -260
rect 7540 -270 7600 -260
rect 7180 -340 7210 -300
rect 7210 -340 7240 -300
rect 7280 -340 7290 -300
rect 7290 -340 7330 -300
rect 7330 -340 7340 -300
rect 7440 -340 7450 -300
rect 7450 -340 7490 -300
rect 7490 -340 7500 -300
rect 7540 -340 7570 -300
rect 7570 -340 7600 -300
rect 7180 -360 7240 -340
rect 7280 -360 7340 -340
rect 7440 -360 7500 -340
rect 7540 -360 7600 -340
rect 1150 -860 1220 -790
rect 1260 -860 1330 -790
rect 1370 -860 1440 -790
rect 1480 -860 1550 -790
rect 1590 -860 1660 -790
rect 1700 -860 1770 -790
rect 1810 -860 1880 -790
rect 1920 -860 1990 -790
rect 2030 -860 2100 -790
rect 2140 -860 2210 -790
rect 2250 -860 2320 -790
rect 2360 -860 2430 -790
rect 2470 -860 2540 -790
rect 2580 -860 2650 -790
rect 1150 -970 1220 -900
rect 1260 -970 1330 -900
rect 1370 -970 1440 -900
rect 1480 -970 1550 -900
rect 1590 -970 1660 -900
rect 1700 -970 1770 -900
rect 1810 -970 1880 -900
rect 1920 -970 1990 -900
rect 2030 -970 2100 -900
rect 2140 -970 2210 -900
rect 2250 -970 2320 -900
rect 2360 -970 2430 -900
rect 2470 -970 2540 -900
rect 2580 -970 2650 -900
rect 20380 -90 20450 -20
rect 20490 -90 20560 -20
rect 20600 -90 20670 -20
rect 20710 -90 20780 -20
rect 14660 -180 14690 -140
rect 14690 -180 14730 -140
rect 14770 -180 14810 -140
rect 14810 -180 14840 -140
rect 14880 -180 14890 -140
rect 14890 -180 14930 -140
rect 14930 -180 14950 -140
rect 14990 -180 15010 -140
rect 15010 -180 15050 -140
rect 15050 -180 15060 -140
rect 14660 -210 14730 -180
rect 14770 -210 14840 -180
rect 14880 -210 14950 -180
rect 14990 -210 15060 -180
rect 20380 -200 20450 -130
rect 20490 -200 20560 -130
rect 20600 -200 20670 -130
rect 20710 -200 20780 -130
rect 14660 -300 14730 -270
rect 14770 -300 14840 -270
rect 14880 -300 14950 -270
rect 14990 -300 15060 -270
rect 14660 -340 14690 -300
rect 14690 -340 14730 -300
rect 14770 -340 14810 -300
rect 14810 -340 14840 -300
rect 14880 -340 14890 -300
rect 14890 -340 14930 -300
rect 14930 -340 14950 -300
rect 14990 -340 15010 -300
rect 15010 -340 15050 -300
rect 15050 -340 15060 -300
rect 20380 -310 20450 -240
rect 20490 -310 20560 -240
rect 20600 -310 20670 -240
rect 20710 -310 20780 -240
rect 12250 -860 12320 -790
rect 12360 -860 12430 -790
rect 12470 -860 12540 -790
rect 12580 -860 12650 -790
rect 12690 -860 12760 -790
rect 12800 -860 12870 -790
rect 12910 -860 12980 -790
rect 13020 -860 13090 -790
rect 13130 -860 13200 -790
rect 13240 -860 13310 -790
rect 13350 -860 13420 -790
rect 13460 -860 13530 -790
rect 13570 -860 13640 -790
rect 13680 -860 13750 -790
rect 12250 -970 12320 -900
rect 12360 -970 12430 -900
rect 12470 -970 12540 -900
rect 12580 -970 12650 -900
rect 12690 -970 12760 -900
rect 12800 -970 12870 -900
rect 12910 -970 12980 -900
rect 13020 -970 13090 -900
rect 13130 -970 13200 -900
rect 13240 -970 13310 -900
rect 13350 -970 13420 -900
rect 13460 -970 13530 -900
rect 13570 -970 13640 -900
rect 13680 -970 13750 -900
rect 25310 -1490 25370 -1430
rect 25410 -1490 25470 -1430
rect 25510 -1490 25570 -1430
rect 25310 -1590 25370 -1530
rect 25410 -1590 25470 -1530
rect 25510 -1590 25570 -1530
rect 25310 -1690 25370 -1630
rect 25410 -1690 25470 -1630
rect 25510 -1690 25570 -1630
rect 25310 -1790 25370 -1730
rect 25410 -1790 25470 -1730
rect 25510 -1790 25570 -1730
rect 25310 -1890 25370 -1830
rect 25410 -1890 25470 -1830
rect 25510 -1890 25570 -1830
rect 25310 -1990 25370 -1930
rect 25410 -1990 25470 -1930
rect 25510 -1990 25570 -1930
rect 25310 -2090 25370 -2030
rect 25410 -2090 25470 -2030
rect 25510 -2090 25570 -2030
rect 25310 -2190 25370 -2130
rect 25410 -2190 25470 -2130
rect 25510 -2190 25570 -2130
rect 25310 -2290 25370 -2230
rect 25410 -2290 25470 -2230
rect 25510 -2290 25570 -2230
rect 1570 -2850 1640 -2780
rect 1680 -2850 1750 -2780
rect 1790 -2850 1860 -2780
rect 1900 -2850 1970 -2780
rect 2010 -2850 2080 -2780
rect 2120 -2850 2190 -2780
rect 2230 -2850 2300 -2780
rect 2340 -2850 2410 -2780
rect 2450 -2850 2520 -2780
rect 2560 -2850 2630 -2780
rect 2670 -2850 2740 -2780
rect 2780 -2850 2850 -2780
rect 2890 -2850 2960 -2780
rect 3000 -2850 3070 -2780
rect 1570 -2960 1640 -2890
rect 1680 -2960 1750 -2890
rect 1790 -2960 1860 -2890
rect 1900 -2960 1970 -2890
rect 2010 -2960 2080 -2890
rect 2120 -2960 2190 -2890
rect 2230 -2960 2300 -2890
rect 2340 -2960 2410 -2890
rect 2450 -2960 2520 -2890
rect 2560 -2960 2630 -2890
rect 2670 -2960 2740 -2890
rect 2780 -2960 2850 -2890
rect 2890 -2960 2960 -2890
rect 3000 -2960 3070 -2890
rect 11790 -2850 11860 -2780
rect 11900 -2850 11970 -2780
rect 12010 -2850 12080 -2780
rect 12120 -2850 12190 -2780
rect 12230 -2850 12300 -2780
rect 12340 -2850 12410 -2780
rect 12450 -2850 12520 -2780
rect 12560 -2850 12630 -2780
rect 12670 -2850 12740 -2780
rect 12780 -2850 12850 -2780
rect 12890 -2850 12960 -2780
rect 13000 -2850 13070 -2780
rect 13110 -2850 13180 -2780
rect 13220 -2850 13290 -2780
rect 11790 -2960 11860 -2890
rect 11900 -2960 11970 -2890
rect 12010 -2960 12080 -2890
rect 12120 -2960 12190 -2890
rect 12230 -2960 12300 -2890
rect 12340 -2960 12410 -2890
rect 12450 -2960 12520 -2890
rect 12560 -2960 12630 -2890
rect 12670 -2960 12740 -2890
rect 12780 -2960 12850 -2890
rect 12890 -2960 12960 -2890
rect 13000 -2960 13070 -2890
rect 13110 -2960 13180 -2890
rect 13220 -2960 13290 -2890
rect 22340 -3120 22410 -3050
rect 22450 -3120 22520 -3050
rect 22560 -3120 22630 -3050
rect 22340 -3230 22410 -3160
rect 22450 -3230 22520 -3160
rect 22560 -3230 22630 -3160
rect 22340 -3340 22410 -3270
rect 22450 -3340 22520 -3270
rect 22560 -3340 22630 -3270
rect 7380 -3400 7440 -3340
rect 7480 -3400 7540 -3340
rect 7380 -3550 7440 -3440
rect 7480 -3550 7540 -3440
rect 7380 -3650 7440 -3590
rect 7480 -3650 7540 -3590
rect 20070 -3760 20140 -3690
rect 20180 -3760 20250 -3690
rect 20290 -3760 20360 -3690
rect 20400 -3760 20470 -3690
rect 20070 -3870 20140 -3800
rect 20180 -3870 20250 -3800
rect 20290 -3870 20360 -3800
rect 20400 -3870 20470 -3800
rect 24550 -3760 24620 -3690
rect 24660 -3760 24730 -3690
rect 24770 -3760 24840 -3690
rect 24880 -3760 24950 -3690
rect 24550 -3870 24620 -3800
rect 24660 -3870 24730 -3800
rect 24770 -3870 24840 -3800
rect 24880 -3870 24950 -3800
rect -2200 -4480 -2178 -4470
rect -2178 -4480 -2138 -4470
rect -2138 -4480 -2130 -4470
rect -2090 -4480 -2058 -4470
rect -2058 -4480 -2020 -4470
rect -2200 -4520 -2130 -4480
rect -2090 -4520 -2020 -4480
rect -2200 -4540 -2178 -4520
rect -2178 -4540 -2138 -4520
rect -2138 -4540 -2130 -4520
rect -2090 -4540 -2058 -4520
rect -2058 -4540 -2020 -4520
rect -2200 -4600 -2130 -4580
rect -2090 -4600 -2020 -4580
rect -2200 -4640 -2178 -4600
rect -2178 -4640 -2138 -4600
rect -2138 -4640 -2130 -4600
rect -2090 -4640 -2058 -4600
rect -2058 -4640 -2020 -4600
rect -2200 -4650 -2130 -4640
rect -2090 -4650 -2020 -4640
rect -2200 -4720 -2178 -4690
rect -2178 -4720 -2138 -4690
rect -2138 -4720 -2130 -4690
rect -2090 -4720 -2058 -4690
rect -2058 -4720 -2020 -4690
rect -2200 -4760 -2130 -4720
rect -2090 -4760 -2020 -4720
rect -2200 -4840 -2130 -4800
rect -2090 -4840 -2020 -4800
rect -2200 -4870 -2178 -4840
rect -2178 -4870 -2138 -4840
rect -2138 -4870 -2130 -4840
rect -2090 -4870 -2058 -4840
rect -2058 -4870 -2020 -4840
rect 7310 -4630 7380 -4560
rect 7420 -4630 7490 -4560
rect 7530 -4630 7600 -4560
rect 7310 -4740 7380 -4670
rect 7420 -4740 7490 -4670
rect 7530 -4740 7600 -4670
rect 7310 -4850 7380 -4780
rect 7420 -4850 7490 -4780
rect 7530 -4850 7600 -4780
rect -2140 -5280 -2070 -5240
rect -2030 -5280 -1960 -5240
rect -2140 -5310 -2138 -5280
rect -2138 -5310 -2098 -5280
rect -2098 -5310 -2070 -5280
rect -2030 -5310 -2018 -5280
rect -2018 -5310 -1978 -5280
rect -1978 -5310 -1960 -5280
rect -2140 -5360 -2070 -5350
rect -2030 -5360 -1960 -5350
rect -2140 -5400 -2138 -5360
rect -2138 -5400 -2098 -5360
rect -2098 -5400 -2070 -5360
rect -2030 -5400 -2018 -5360
rect -2018 -5400 -1978 -5360
rect -1978 -5400 -1960 -5360
rect -2140 -5420 -2070 -5400
rect -2030 -5420 -1960 -5400
rect -2140 -5480 -2138 -5460
rect -2138 -5480 -2098 -5460
rect -2098 -5480 -2070 -5460
rect -2030 -5480 -2018 -5460
rect -2018 -5480 -1978 -5460
rect -1978 -5480 -1960 -5460
rect -2140 -5520 -2070 -5480
rect -2030 -5520 -1960 -5480
rect -2140 -5530 -2138 -5520
rect -2138 -5530 -2098 -5520
rect -2098 -5530 -2070 -5520
rect -2030 -5530 -2018 -5520
rect -2018 -5530 -1978 -5520
rect -1978 -5530 -1960 -5520
rect -2140 -5600 -2070 -5570
rect -2030 -5600 -1960 -5570
rect -2140 -5640 -2138 -5600
rect -2138 -5640 -2098 -5600
rect -2098 -5640 -2070 -5600
rect -2030 -5640 -2018 -5600
rect -2018 -5640 -1978 -5600
rect -1978 -5640 -1960 -5600
rect -840 -6530 -800 -6500
rect -800 -6530 -770 -6500
rect -710 -6530 -680 -6500
rect -680 -6530 -640 -6500
rect -840 -6570 -770 -6530
rect -710 -6570 -640 -6530
rect -840 -6650 -770 -6610
rect -710 -6650 -640 -6610
rect -840 -6680 -800 -6650
rect -800 -6680 -770 -6650
rect -710 -6680 -680 -6650
rect -680 -6680 -640 -6650
rect 7050 -6520 7110 -6460
rect 7150 -6520 7210 -6460
rect 7250 -6520 7310 -6460
rect 7590 -6520 7650 -6460
rect 7690 -6520 7750 -6460
rect 7790 -6520 7850 -6460
rect 7050 -6620 7110 -6560
rect 7150 -6620 7210 -6560
rect 7250 -6620 7310 -6560
rect 7590 -6620 7650 -6560
rect 7690 -6620 7750 -6560
rect 7790 -6620 7850 -6560
rect -840 -6730 -770 -6720
rect -710 -6730 -640 -6720
rect -840 -6770 -800 -6730
rect -800 -6770 -770 -6730
rect -710 -6770 -680 -6730
rect -680 -6770 -640 -6730
rect -840 -6790 -770 -6770
rect -710 -6790 -640 -6770
rect 4770 -6730 4830 -6670
rect 4870 -6730 4930 -6670
rect 4970 -6730 5030 -6670
rect 7050 -6720 7110 -6660
rect 7150 -6720 7210 -6660
rect 7250 -6720 7310 -6660
rect 7590 -6720 7650 -6660
rect 7690 -6720 7750 -6660
rect 7790 -6720 7850 -6660
rect 9870 -6730 9930 -6670
rect 9970 -6730 10030 -6670
rect 10070 -6730 10130 -6670
rect 15420 -6530 15460 -6500
rect 15460 -6530 15490 -6500
rect 15550 -6530 15580 -6500
rect 15580 -6530 15620 -6500
rect 15420 -6570 15490 -6530
rect 15550 -6570 15620 -6530
rect 15420 -6650 15490 -6610
rect 15550 -6650 15620 -6610
rect 15420 -6680 15460 -6650
rect 15460 -6680 15490 -6650
rect 15550 -6680 15580 -6650
rect 15580 -6680 15620 -6650
rect -840 -6850 -800 -6830
rect -800 -6850 -770 -6830
rect -710 -6850 -680 -6830
rect -680 -6850 -640 -6830
rect -840 -6890 -770 -6850
rect -710 -6890 -640 -6850
rect -840 -6900 -800 -6890
rect -800 -6900 -770 -6890
rect -710 -6900 -680 -6890
rect -680 -6900 -640 -6890
rect 4770 -6830 4830 -6770
rect 4870 -6830 4930 -6770
rect 4970 -6830 5030 -6770
rect 7050 -6820 7110 -6760
rect 7150 -6820 7210 -6760
rect 7250 -6820 7310 -6760
rect 7590 -6820 7650 -6760
rect 7690 -6820 7750 -6760
rect 7790 -6820 7850 -6760
rect 9870 -6830 9930 -6770
rect 9970 -6830 10030 -6770
rect 10070 -6830 10130 -6770
rect 15420 -6730 15490 -6720
rect 15550 -6730 15620 -6720
rect 15420 -6770 15460 -6730
rect 15460 -6770 15490 -6730
rect 15550 -6770 15580 -6730
rect 15580 -6770 15620 -6730
rect 15420 -6790 15490 -6770
rect 15550 -6790 15620 -6770
rect 4770 -6930 4830 -6870
rect 4870 -6930 4930 -6870
rect 4970 -6930 5030 -6870
rect 9870 -6930 9930 -6870
rect 9970 -6930 10030 -6870
rect 10070 -6930 10130 -6870
rect 15420 -6850 15460 -6830
rect 15460 -6850 15490 -6830
rect 15550 -6850 15580 -6830
rect 15580 -6850 15620 -6830
rect 15420 -6890 15490 -6850
rect 15550 -6890 15620 -6850
rect 15420 -6900 15460 -6890
rect 15460 -6900 15490 -6890
rect 15550 -6900 15580 -6890
rect 15580 -6900 15620 -6890
rect -2200 -7880 -2178 -7870
rect -2178 -7880 -2138 -7870
rect -2138 -7880 -2130 -7870
rect -2090 -7880 -2058 -7870
rect -2058 -7880 -2020 -7870
rect -2200 -7920 -2130 -7880
rect -2090 -7920 -2020 -7880
rect -2200 -7940 -2178 -7920
rect -2178 -7940 -2138 -7920
rect -2138 -7940 -2130 -7920
rect -2090 -7940 -2058 -7920
rect -2058 -7940 -2020 -7920
rect -2200 -8000 -2130 -7980
rect -2090 -8000 -2020 -7980
rect -2200 -8040 -2178 -8000
rect -2178 -8040 -2138 -8000
rect -2138 -8040 -2130 -8000
rect -2090 -8040 -2058 -8000
rect -2058 -8040 -2020 -8000
rect -2200 -8050 -2130 -8040
rect -2090 -8050 -2020 -8040
rect -2200 -8120 -2178 -8090
rect -2178 -8120 -2138 -8090
rect -2138 -8120 -2130 -8090
rect -2090 -8120 -2058 -8090
rect -2058 -8120 -2020 -8090
rect -2200 -8160 -2130 -8120
rect -2090 -8160 -2020 -8120
rect -2200 -8240 -2130 -8200
rect -2090 -8240 -2020 -8200
rect -2200 -8270 -2178 -8240
rect -2178 -8270 -2138 -8240
rect -2138 -8270 -2130 -8240
rect -2090 -8270 -2058 -8240
rect -2058 -8270 -2020 -8240
rect 14600 -8300 14670 -8230
rect 14700 -8300 14770 -8230
rect 14810 -8300 14880 -8230
rect 14600 -8410 14670 -8340
rect 14700 -8410 14770 -8340
rect 14810 -8410 14880 -8340
rect 14600 -8520 14670 -8450
rect 14700 -8520 14770 -8450
rect 14810 -8520 14880 -8450
rect -2140 -8680 -2070 -8640
rect -2030 -8680 -1960 -8640
rect -2140 -8710 -2138 -8680
rect -2138 -8710 -2098 -8680
rect -2098 -8710 -2070 -8680
rect -2030 -8710 -2018 -8680
rect -2018 -8710 -1978 -8680
rect -1978 -8710 -1960 -8680
rect -2140 -8760 -2070 -8750
rect -2030 -8760 -1960 -8750
rect -2140 -8800 -2138 -8760
rect -2138 -8800 -2098 -8760
rect -2098 -8800 -2070 -8760
rect -2030 -8800 -2018 -8760
rect -2018 -8800 -1978 -8760
rect -1978 -8800 -1960 -8760
rect -2140 -8820 -2070 -8800
rect -2030 -8820 -1960 -8800
rect 19230 -8630 19300 -8560
rect 19330 -8630 19400 -8560
rect 19430 -8630 19500 -8560
rect 19230 -8730 19300 -8660
rect 19330 -8730 19400 -8660
rect 19430 -8730 19500 -8660
rect 19230 -8830 19300 -8760
rect 19330 -8830 19400 -8760
rect 19430 -8830 19500 -8760
rect -2140 -8880 -2138 -8860
rect -2138 -8880 -2098 -8860
rect -2098 -8880 -2070 -8860
rect -2030 -8880 -2018 -8860
rect -2018 -8880 -1978 -8860
rect -1978 -8880 -1960 -8860
rect -2140 -8920 -2070 -8880
rect -2030 -8920 -1960 -8880
rect -2140 -8930 -2138 -8920
rect -2138 -8930 -2098 -8920
rect -2098 -8930 -2070 -8920
rect -2030 -8930 -2018 -8920
rect -2018 -8930 -1978 -8920
rect -1978 -8930 -1960 -8920
rect -2140 -9000 -2070 -8970
rect -2030 -9000 -1960 -8970
rect -2140 -9040 -2138 -9000
rect -2138 -9040 -2098 -9000
rect -2098 -9040 -2070 -9000
rect -2030 -9040 -2018 -9000
rect -2018 -9040 -1978 -9000
rect -1978 -9040 -1960 -9000
rect 19960 -9070 20030 -9000
rect 20060 -9070 20130 -9000
rect 20160 -9070 20230 -9000
rect 19960 -9170 20030 -9100
rect 20060 -9170 20130 -9100
rect 20160 -9170 20230 -9100
rect 19960 -9270 20030 -9200
rect 20060 -9270 20130 -9200
rect 20160 -9270 20230 -9200
rect -240 -9700 -210 -9660
rect -210 -9700 -170 -9660
rect -130 -9700 -90 -9660
rect -90 -9700 -60 -9660
rect -20 -9700 -10 -9660
rect -10 -9700 30 -9660
rect 30 -9700 50 -9660
rect 90 -9700 110 -9660
rect 110 -9700 150 -9660
rect 150 -9700 160 -9660
rect -240 -9730 -170 -9700
rect -130 -9730 -60 -9700
rect -20 -9730 50 -9700
rect 90 -9730 160 -9700
rect -240 -9820 -170 -9790
rect -130 -9820 -60 -9790
rect -20 -9820 50 -9790
rect 90 -9820 160 -9790
rect -240 -9860 -210 -9820
rect -210 -9860 -170 -9820
rect -130 -9860 -90 -9820
rect -90 -9860 -60 -9820
rect -20 -9860 -10 -9820
rect -10 -9860 30 -9820
rect 30 -9860 50 -9820
rect 90 -9860 110 -9820
rect 110 -9860 150 -9820
rect 150 -9860 160 -9820
rect 7240 -9660 7300 -9640
rect 7340 -9660 7400 -9640
rect 7500 -9660 7560 -9640
rect 7600 -9660 7660 -9640
rect 7240 -9700 7270 -9660
rect 7270 -9700 7300 -9660
rect 7340 -9700 7350 -9660
rect 7350 -9700 7390 -9660
rect 7390 -9700 7400 -9660
rect 7500 -9700 7510 -9660
rect 7510 -9700 7550 -9660
rect 7550 -9700 7560 -9660
rect 7600 -9700 7630 -9660
rect 7630 -9700 7660 -9660
rect 7240 -9740 7300 -9730
rect 7340 -9740 7400 -9730
rect 7500 -9740 7560 -9730
rect 7600 -9740 7660 -9730
rect 7240 -9780 7270 -9740
rect 7270 -9780 7300 -9740
rect 7340 -9780 7350 -9740
rect 7350 -9780 7390 -9740
rect 7390 -9780 7400 -9740
rect 7500 -9780 7510 -9740
rect 7510 -9780 7550 -9740
rect 7550 -9780 7560 -9740
rect 7600 -9780 7630 -9740
rect 7630 -9780 7660 -9740
rect 7240 -9790 7300 -9780
rect 7340 -9790 7400 -9780
rect 7500 -9790 7560 -9780
rect 7600 -9790 7660 -9780
rect 7240 -9860 7270 -9820
rect 7270 -9860 7300 -9820
rect 7340 -9860 7350 -9820
rect 7350 -9860 7390 -9820
rect 7390 -9860 7400 -9820
rect 7500 -9860 7510 -9820
rect 7510 -9860 7550 -9820
rect 7550 -9860 7560 -9820
rect 7600 -9860 7630 -9820
rect 7630 -9860 7660 -9820
rect 7240 -9880 7300 -9860
rect 7340 -9880 7400 -9860
rect 7500 -9880 7560 -9860
rect 7600 -9880 7660 -9860
rect 1150 -10410 1220 -10340
rect 1260 -10410 1330 -10340
rect 1370 -10410 1440 -10340
rect 1480 -10410 1550 -10340
rect 1590 -10410 1660 -10340
rect 1700 -10410 1770 -10340
rect 1810 -10410 1880 -10340
rect 1920 -10410 1990 -10340
rect 2030 -10410 2100 -10340
rect 2140 -10410 2210 -10340
rect 2250 -10410 2320 -10340
rect 2360 -10410 2430 -10340
rect 2470 -10410 2540 -10340
rect 2580 -10410 2650 -10340
rect 1150 -10520 1220 -10450
rect 1260 -10520 1330 -10450
rect 1370 -10520 1440 -10450
rect 1480 -10520 1550 -10450
rect 1590 -10520 1660 -10450
rect 1700 -10520 1770 -10450
rect 1810 -10520 1880 -10450
rect 1920 -10520 1990 -10450
rect 2030 -10520 2100 -10450
rect 2140 -10520 2210 -10450
rect 2250 -10520 2320 -10450
rect 2360 -10520 2430 -10450
rect 2470 -10520 2540 -10450
rect 2580 -10520 2650 -10450
rect 14720 -9700 14750 -9660
rect 14750 -9700 14790 -9660
rect 14830 -9700 14870 -9660
rect 14870 -9700 14900 -9660
rect 14940 -9700 14950 -9660
rect 14950 -9700 14990 -9660
rect 14990 -9700 15010 -9660
rect 15050 -9700 15070 -9660
rect 15070 -9700 15110 -9660
rect 15110 -9700 15120 -9660
rect 14720 -9730 14790 -9700
rect 14830 -9730 14900 -9700
rect 14940 -9730 15010 -9700
rect 15050 -9730 15120 -9700
rect 14720 -9820 14790 -9790
rect 14830 -9820 14900 -9790
rect 14940 -9820 15010 -9790
rect 15050 -9820 15120 -9790
rect 14720 -9860 14750 -9820
rect 14750 -9860 14790 -9820
rect 14830 -9860 14870 -9820
rect 14870 -9860 14900 -9820
rect 14940 -9860 14950 -9820
rect 14950 -9860 14990 -9820
rect 14990 -9860 15010 -9820
rect 15050 -9860 15070 -9820
rect 15070 -9860 15110 -9820
rect 15110 -9860 15120 -9820
rect 12290 -10440 12360 -10370
rect 12400 -10440 12470 -10370
rect 12510 -10440 12580 -10370
rect 12620 -10440 12690 -10370
rect 12730 -10440 12800 -10370
rect 12840 -10440 12910 -10370
rect 12950 -10440 13020 -10370
rect 13060 -10440 13130 -10370
rect 13170 -10440 13240 -10370
rect 13280 -10440 13350 -10370
rect 13390 -10440 13460 -10370
rect 13500 -10440 13570 -10370
rect 13610 -10440 13680 -10370
rect 13720 -10440 13790 -10370
rect 12290 -10550 12360 -10480
rect 12400 -10550 12470 -10480
rect 12510 -10550 12580 -10480
rect 12620 -10550 12690 -10480
rect 12730 -10550 12800 -10480
rect 12840 -10550 12910 -10480
rect 12950 -10550 13020 -10480
rect 13060 -10550 13130 -10480
rect 13170 -10550 13240 -10480
rect 13280 -10550 13350 -10480
rect 13390 -10550 13460 -10480
rect 13500 -10550 13570 -10480
rect 13610 -10550 13680 -10480
rect 13720 -10550 13790 -10480
rect 2240 -12370 2310 -12300
rect 2350 -12370 2420 -12300
rect 2460 -12370 2530 -12300
rect 2570 -12370 2640 -12300
rect 2680 -12370 2750 -12300
rect 2790 -12370 2860 -12300
rect 2900 -12370 2970 -12300
rect 3010 -12370 3080 -12300
rect 3120 -12370 3190 -12300
rect 3230 -12370 3300 -12300
rect 3340 -12370 3410 -12300
rect 3450 -12370 3520 -12300
rect 3560 -12370 3630 -12300
rect 3670 -12370 3740 -12300
rect 2240 -12480 2310 -12410
rect 2350 -12480 2420 -12410
rect 2460 -12480 2530 -12410
rect 2570 -12480 2640 -12410
rect 2680 -12480 2750 -12410
rect 2790 -12480 2860 -12410
rect 2900 -12480 2970 -12410
rect 3010 -12480 3080 -12410
rect 3120 -12480 3190 -12410
rect 3230 -12480 3300 -12410
rect 3340 -12480 3410 -12410
rect 3450 -12480 3520 -12410
rect 3560 -12480 3630 -12410
rect 3670 -12480 3740 -12410
rect 11120 -12370 11190 -12300
rect 11230 -12370 11300 -12300
rect 11340 -12370 11410 -12300
rect 11450 -12370 11520 -12300
rect 11560 -12370 11630 -12300
rect 11670 -12370 11740 -12300
rect 11780 -12370 11850 -12300
rect 11890 -12370 11960 -12300
rect 12000 -12370 12070 -12300
rect 12110 -12370 12180 -12300
rect 12220 -12370 12290 -12300
rect 12330 -12370 12400 -12300
rect 12440 -12370 12510 -12300
rect 12550 -12370 12620 -12300
rect 11120 -12480 11190 -12410
rect 11230 -12480 11300 -12410
rect 11340 -12480 11410 -12410
rect 11450 -12480 11520 -12410
rect 11560 -12480 11630 -12410
rect 11670 -12480 11740 -12410
rect 11780 -12480 11850 -12410
rect 11890 -12480 11960 -12410
rect 12000 -12480 12070 -12410
rect 12110 -12480 12180 -12410
rect 12220 -12480 12290 -12410
rect 12330 -12480 12400 -12410
rect 12440 -12480 12510 -12410
rect 12550 -12480 12620 -12410
rect 7010 -13310 7070 -13250
rect 7110 -13310 7170 -13250
rect 7210 -13310 7270 -13250
rect 7630 -13310 7690 -13250
rect 7730 -13310 7790 -13250
rect 7830 -13310 7890 -13250
rect 7010 -13400 7070 -13340
rect 7110 -13400 7170 -13340
rect 7210 -13400 7270 -13340
rect 7630 -13400 7690 -13340
rect 7730 -13400 7790 -13340
rect 7830 -13400 7890 -13340
rect 7010 -13490 7070 -13430
rect 7110 -13490 7170 -13430
rect 7210 -13490 7270 -13430
rect 7630 -13490 7690 -13430
rect 7730 -13490 7790 -13430
rect 7830 -13490 7890 -13430
rect 7010 -13590 7070 -13530
rect 7110 -13590 7170 -13530
rect 7210 -13590 7270 -13530
rect 7630 -13590 7690 -13530
rect 7730 -13590 7790 -13530
rect 7830 -13590 7890 -13530
rect 7010 -13680 7070 -13620
rect 7110 -13680 7170 -13620
rect 7210 -13680 7270 -13620
rect 7630 -13680 7690 -13620
rect 7730 -13680 7790 -13620
rect 7830 -13680 7890 -13620
rect 7010 -13770 7070 -13710
rect 7110 -13770 7170 -13710
rect 7210 -13770 7270 -13710
rect 7630 -13770 7690 -13710
rect 7730 -13770 7790 -13710
rect 7830 -13770 7890 -13710
rect 19230 -14290 19300 -14220
rect 19330 -14290 19400 -14220
rect 19430 -14290 19500 -14220
rect 19230 -14390 19300 -14320
rect 19330 -14390 19400 -14320
rect 19430 -14390 19500 -14320
rect 19230 -14490 19300 -14420
rect 19330 -14490 19400 -14420
rect 19430 -14490 19500 -14420
rect 20480 -14940 20550 -14870
rect 20580 -14940 20650 -14870
rect 20680 -14940 20750 -14870
rect 20480 -15040 20550 -14970
rect 20580 -15040 20650 -14970
rect 20680 -15040 20750 -14970
rect 20480 -15140 20550 -15070
rect 20580 -15140 20650 -15070
rect 20680 -15140 20750 -15070
rect 5040 -17160 5100 -17100
rect 5140 -17160 5200 -17100
rect 5240 -17160 5300 -17100
rect 9600 -17160 9660 -17100
rect 9700 -17160 9760 -17100
rect 9800 -17160 9860 -17100
rect 5040 -17260 5100 -17200
rect 5140 -17260 5200 -17200
rect 5240 -17260 5300 -17200
rect 9600 -17260 9660 -17200
rect 9700 -17260 9760 -17200
rect 9800 -17260 9860 -17200
rect 5040 -17360 5100 -17300
rect 5140 -17360 5200 -17300
rect 5240 -17360 5300 -17300
rect 9600 -17360 9660 -17300
rect 9700 -17360 9760 -17300
rect 9800 -17360 9860 -17300
rect 7230 -17670 7300 -17600
rect 7340 -17670 7410 -17600
rect 7450 -17670 7520 -17600
rect 7560 -17670 7630 -17600
rect 7230 -17780 7300 -17710
rect 7340 -17780 7410 -17710
rect 7450 -17780 7520 -17710
rect 7560 -17780 7630 -17710
rect 7230 -17890 7300 -17820
rect 7340 -17890 7410 -17820
rect 7450 -17890 7520 -17820
rect 7560 -17890 7630 -17820
rect 7230 -18000 7300 -17930
rect 7340 -18000 7410 -17930
rect 7450 -18000 7520 -17930
rect 7560 -18000 7630 -17930
rect 19230 -20360 19300 -20290
rect 19330 -20360 19400 -20290
rect 19430 -20360 19500 -20290
rect 19230 -20460 19300 -20390
rect 19330 -20460 19400 -20390
rect 19430 -20460 19500 -20390
rect 19230 -20560 19300 -20490
rect 19330 -20560 19400 -20490
rect 19430 -20560 19500 -20490
rect 20040 -20790 20110 -20720
rect 20140 -20790 20210 -20720
rect 20240 -20790 20310 -20720
rect 20040 -20890 20110 -20820
rect 20140 -20890 20210 -20820
rect 20240 -20890 20310 -20820
rect 20040 -20990 20110 -20920
rect 20140 -20990 20210 -20920
rect 20240 -20990 20310 -20920
rect 2280 -22730 2350 -22660
rect 2390 -22730 2460 -22660
rect 2500 -22730 2570 -22660
rect 2610 -22730 2680 -22660
rect 2720 -22730 2790 -22660
rect 2830 -22730 2900 -22660
rect 2940 -22730 3010 -22660
rect 3050 -22730 3120 -22660
rect 3160 -22730 3230 -22660
rect 3270 -22730 3340 -22660
rect 3380 -22730 3450 -22660
rect 3490 -22730 3560 -22660
rect 3600 -22730 3670 -22660
rect 3710 -22730 3780 -22660
rect 2280 -22840 2350 -22770
rect 2390 -22840 2460 -22770
rect 2500 -22840 2570 -22770
rect 2610 -22840 2680 -22770
rect 2720 -22840 2790 -22770
rect 2830 -22840 2900 -22770
rect 2940 -22840 3010 -22770
rect 3050 -22840 3120 -22770
rect 3160 -22840 3230 -22770
rect 3270 -22840 3340 -22770
rect 3380 -22840 3450 -22770
rect 3490 -22840 3560 -22770
rect 3600 -22840 3670 -22770
rect 3710 -22840 3780 -22770
rect 11160 -22730 11230 -22660
rect 11270 -22730 11340 -22660
rect 11380 -22730 11450 -22660
rect 11490 -22730 11560 -22660
rect 11600 -22730 11670 -22660
rect 11710 -22730 11780 -22660
rect 11820 -22730 11890 -22660
rect 11930 -22730 12000 -22660
rect 12040 -22730 12110 -22660
rect 12150 -22730 12220 -22660
rect 12260 -22730 12330 -22660
rect 12370 -22730 12440 -22660
rect 12480 -22730 12550 -22660
rect 12590 -22730 12660 -22660
rect 11160 -22840 11230 -22770
rect 11270 -22840 11340 -22770
rect 11380 -22840 11450 -22770
rect 11490 -22840 11560 -22770
rect 11600 -22840 11670 -22770
rect 11710 -22840 11780 -22770
rect 11820 -22840 11890 -22770
rect 11930 -22840 12000 -22770
rect 12040 -22840 12110 -22770
rect 12150 -22840 12220 -22770
rect 12260 -22840 12330 -22770
rect 12370 -22840 12440 -22770
rect 12480 -22840 12550 -22770
rect 12590 -22840 12660 -22770
<< metal2 >>
rect 21060 7210 21540 7260
rect 21060 7140 21090 7210
rect 21160 7140 21200 7210
rect 21270 7140 21310 7210
rect 21380 7140 21420 7210
rect 21490 7140 21540 7210
rect 21060 7100 21540 7140
rect 21060 7030 21090 7100
rect 21160 7030 21200 7100
rect 21270 7030 21310 7100
rect 21380 7030 21420 7100
rect 21490 7030 21540 7100
rect 21060 7000 21540 7030
rect 23460 7210 23940 7260
rect 23460 7140 23490 7210
rect 23560 7140 23600 7210
rect 23670 7140 23710 7210
rect 23780 7140 23820 7210
rect 23890 7140 23940 7210
rect 23460 7100 23940 7140
rect 23460 7030 23490 7100
rect 23560 7030 23600 7100
rect 23670 7030 23710 7100
rect 23780 7030 23820 7100
rect 23890 7030 23940 7100
rect 23460 7000 23940 7030
rect 1540 6850 3140 6900
rect 1540 6780 1570 6850
rect 1640 6780 1680 6850
rect 1750 6780 1790 6850
rect 1860 6780 1900 6850
rect 1970 6780 2010 6850
rect 2080 6780 2120 6850
rect 2190 6780 2230 6850
rect 2300 6780 2340 6850
rect 2410 6780 2450 6850
rect 2520 6780 2560 6850
rect 2630 6780 2670 6850
rect 2740 6780 2780 6850
rect 2850 6780 2890 6850
rect 2960 6780 3000 6850
rect 3070 6780 3140 6850
rect 1540 6740 3140 6780
rect 1540 6670 1570 6740
rect 1640 6670 1680 6740
rect 1750 6670 1790 6740
rect 1860 6670 1900 6740
rect 1970 6670 2010 6740
rect 2080 6670 2120 6740
rect 2190 6670 2230 6740
rect 2300 6670 2340 6740
rect 2410 6670 2450 6740
rect 2520 6670 2560 6740
rect 2630 6670 2670 6740
rect 2740 6670 2780 6740
rect 2850 6670 2890 6740
rect 2960 6670 3000 6740
rect 3070 6670 3140 6740
rect 11760 6880 13360 6930
rect 11760 6810 11790 6880
rect 11860 6810 11900 6880
rect 11970 6810 12010 6880
rect 12080 6810 12120 6880
rect 12190 6810 12230 6880
rect 12300 6810 12340 6880
rect 12410 6810 12450 6880
rect 12520 6810 12560 6880
rect 12630 6810 12670 6880
rect 12740 6810 12780 6880
rect 12850 6810 12890 6880
rect 12960 6810 13000 6880
rect 13070 6810 13110 6880
rect 13180 6810 13220 6880
rect 13290 6810 13360 6880
rect 11760 6770 13360 6810
rect 11760 6700 11790 6770
rect 11860 6700 11900 6770
rect 11970 6700 12010 6770
rect 12080 6700 12120 6770
rect 12190 6700 12230 6770
rect 12300 6700 12340 6770
rect 12410 6700 12450 6770
rect 12520 6700 12560 6770
rect 12630 6700 12670 6770
rect 12740 6700 12780 6770
rect 12850 6700 12890 6770
rect 12960 6700 13000 6770
rect 13070 6700 13110 6770
rect 13180 6700 13220 6770
rect 13290 6700 13360 6770
rect 11760 6670 13360 6700
rect 1540 6640 3140 6670
rect 7350 6300 28540 6320
rect 7350 6290 28340 6300
rect 7350 6230 7380 6290
rect 7440 6230 7480 6290
rect 7540 6280 28340 6290
rect 7540 6230 20380 6280
rect 7350 6210 20380 6230
rect 20450 6210 20490 6280
rect 20560 6210 20600 6280
rect 20670 6210 20710 6280
rect 20780 6230 28340 6280
rect 28410 6230 28450 6300
rect 28520 6230 28540 6300
rect 20780 6210 28540 6230
rect 7350 6190 28540 6210
rect 7350 6080 7380 6190
rect 7440 6080 7480 6190
rect 7540 6170 28540 6190
rect 7540 6100 20380 6170
rect 20450 6100 20490 6170
rect 20560 6100 20600 6170
rect 20670 6100 20710 6170
rect 20780 6100 28340 6170
rect 28410 6100 28450 6170
rect 28520 6100 28540 6170
rect 7540 6080 28540 6100
rect 7350 6060 28540 6080
rect 7350 6040 20380 6060
rect 7350 5980 7380 6040
rect 7440 5980 7480 6040
rect 7540 5990 20380 6040
rect 20450 5990 20490 6060
rect 20560 5990 20600 6060
rect 20670 5990 20710 6060
rect 20780 6040 28540 6060
rect 20780 5990 28340 6040
rect 7540 5980 28340 5990
rect 7350 5970 28340 5980
rect 28410 5970 28450 6040
rect 28520 5970 28540 6040
rect 7350 5950 28540 5970
rect 7400 5390 7490 5410
rect 7400 5320 7410 5390
rect 7480 5320 7490 5390
rect 7400 5280 7490 5320
rect 7400 5210 7410 5280
rect 7480 5210 7490 5280
rect 7400 5170 7490 5210
rect 7400 5100 7410 5170
rect 7480 5100 7490 5170
rect 7400 5060 7490 5100
rect 7400 4990 7410 5060
rect 7480 4990 7490 5060
rect 7400 4950 7490 4990
rect 7400 4880 7410 4950
rect 7480 4880 7490 4950
rect 7400 4860 7490 4880
rect 25280 4870 25880 4900
rect 25280 4810 25310 4870
rect 25370 4810 25410 4870
rect 25470 4810 25510 4870
rect 25570 4810 25880 4870
rect 7560 4760 7880 4790
rect 7560 4700 7590 4760
rect 7650 4700 7690 4760
rect 7750 4700 7790 4760
rect 7850 4700 7880 4760
rect 7560 4610 7880 4700
rect 25280 4770 25880 4810
rect 25280 4710 25310 4770
rect 25370 4710 25410 4770
rect 25470 4710 25510 4770
rect 25570 4710 25880 4770
rect 25280 4670 25880 4710
rect 25280 4610 25310 4670
rect 25370 4610 25410 4670
rect 25470 4610 25510 4670
rect 25570 4610 25880 4670
rect -880 4580 -600 4610
rect -880 4510 -840 4580
rect -770 4510 -710 4580
rect -640 4510 -600 4580
rect -880 4470 -600 4510
rect -880 4400 -840 4470
rect -770 4400 -710 4470
rect -640 4400 -600 4470
rect -880 4360 -600 4400
rect -880 4290 -840 4360
rect -770 4290 -710 4360
rect -640 4290 -600 4360
rect -880 4250 -600 4290
rect -880 4180 -840 4250
rect -770 4180 -710 4250
rect -640 4180 -600 4250
rect -880 4130 -600 4180
rect 6670 4580 7880 4610
rect 6670 4520 6700 4580
rect 6760 4520 7880 4580
rect 6670 4460 7880 4520
rect 6670 4400 6700 4460
rect 6760 4400 7880 4460
rect 6670 4340 7880 4400
rect 6670 4280 6700 4340
rect 6760 4280 7880 4340
rect 6670 4220 7880 4280
rect 6670 4160 6700 4220
rect 6760 4160 7880 4220
rect 6670 4130 7880 4160
rect 15380 4580 15660 4610
rect 15380 4510 15420 4580
rect 15490 4510 15550 4580
rect 15620 4510 15660 4580
rect 15380 4470 15660 4510
rect 15380 4400 15420 4470
rect 15490 4400 15550 4470
rect 15620 4400 15660 4470
rect 15380 4360 15660 4400
rect 15380 4290 15420 4360
rect 15490 4290 15550 4360
rect 15620 4290 15660 4360
rect 15380 4250 15660 4290
rect 15380 4180 15420 4250
rect 15490 4180 15550 4250
rect 15620 4180 15660 4250
rect 15380 4130 15660 4180
rect 25280 4570 25880 4610
rect 25280 4510 25310 4570
rect 25370 4510 25410 4570
rect 25470 4510 25510 4570
rect 25570 4510 25880 4570
rect 25280 4470 25880 4510
rect 25280 4410 25310 4470
rect 25370 4410 25410 4470
rect 25470 4410 25510 4470
rect 25570 4410 25880 4470
rect 25280 4370 25880 4410
rect 25280 4310 25310 4370
rect 25370 4310 25410 4370
rect 25470 4310 25510 4370
rect 25570 4310 25880 4370
rect 25280 4270 25880 4310
rect 25280 4210 25310 4270
rect 25370 4210 25410 4270
rect 25470 4210 25510 4270
rect 25570 4210 25880 4270
rect 25280 4170 25880 4210
rect 7020 3240 7340 3270
rect 7020 3180 7050 3240
rect 7110 3180 7150 3240
rect 7210 3180 7250 3240
rect 7310 3180 7340 3240
rect 7020 3140 7340 3180
rect 7020 3080 7050 3140
rect 7110 3080 7150 3140
rect 7210 3080 7250 3140
rect 7310 3080 7340 3140
rect 7020 3040 7340 3080
rect 7020 2980 7050 3040
rect 7110 2980 7150 3040
rect 7210 2980 7250 3040
rect 7310 2980 7340 3040
rect 7020 2960 7340 2980
rect 7560 3240 7880 4130
rect 25280 4110 25310 4170
rect 25370 4110 25410 4170
rect 25470 4110 25510 4170
rect 25570 4110 25880 4170
rect 25280 4070 25880 4110
rect 25280 4010 25310 4070
rect 25370 4010 25410 4070
rect 25470 4010 25510 4070
rect 25570 4010 25880 4070
rect 25280 3980 25880 4010
rect 7560 3180 7590 3240
rect 7650 3180 7690 3240
rect 7750 3180 7790 3240
rect 7850 3180 7880 3240
rect 7560 3140 7880 3180
rect 7560 3080 7590 3140
rect 7650 3080 7690 3140
rect 7750 3080 7790 3140
rect 7850 3080 7880 3140
rect 7560 3040 7880 3080
rect 22300 3360 22630 3380
rect 22300 3290 22320 3360
rect 22390 3290 22430 3360
rect 22500 3290 22540 3360
rect 22610 3290 22630 3360
rect 22300 3250 22630 3290
rect 22300 3180 22320 3250
rect 22390 3180 22430 3250
rect 22500 3180 22540 3250
rect 22610 3180 22630 3250
rect 22300 3140 22630 3180
rect 22300 3070 22320 3140
rect 22390 3070 22430 3140
rect 22500 3070 22540 3140
rect 22610 3070 22630 3140
rect 22300 3050 22630 3070
rect 7560 2980 7590 3040
rect 7650 2980 7690 3040
rect 7750 2980 7790 3040
rect 7850 2980 7880 3040
rect 7560 2960 7880 2980
rect 4740 2890 5060 2920
rect 4740 2830 4770 2890
rect 4830 2830 4870 2890
rect 4930 2830 4970 2890
rect 5030 2830 5060 2890
rect 4740 2790 5060 2830
rect 4740 2730 4770 2790
rect 4830 2730 4870 2790
rect 4930 2730 4970 2790
rect 5030 2730 5060 2790
rect 4740 2690 5060 2730
rect 4740 2630 4770 2690
rect 4830 2630 4870 2690
rect 4930 2630 4970 2690
rect 5030 2630 5060 2690
rect 4740 2610 5060 2630
rect 9840 2890 10160 2920
rect 9840 2830 9870 2890
rect 9930 2830 9970 2890
rect 10030 2830 10070 2890
rect 10130 2830 10160 2890
rect 9840 2790 10160 2830
rect 9840 2730 9870 2790
rect 9930 2730 9970 2790
rect 10030 2730 10070 2790
rect 10130 2730 10160 2790
rect 9840 2690 10160 2730
rect 9840 2630 9870 2690
rect 9930 2630 9970 2690
rect 10030 2630 10070 2690
rect 10130 2630 10160 2690
rect 9840 2610 10160 2630
rect 20020 2600 20500 2630
rect 20020 2530 20070 2600
rect 20140 2530 20180 2600
rect 20250 2530 20290 2600
rect 20360 2530 20400 2600
rect 20470 2530 20500 2600
rect 20020 2490 20500 2530
rect 20020 2420 20070 2490
rect 20140 2420 20180 2490
rect 20250 2420 20290 2490
rect 20360 2420 20400 2490
rect 20470 2420 20500 2490
rect 20020 2370 20500 2420
rect 24500 2600 24980 2630
rect 24500 2530 24550 2600
rect 24620 2530 24660 2600
rect 24730 2530 24770 2600
rect 24840 2530 24880 2600
rect 24950 2530 24980 2600
rect 24500 2490 24980 2530
rect 24500 2420 24550 2490
rect 24620 2420 24660 2490
rect 24730 2420 24770 2490
rect 24840 2420 24880 2490
rect 24950 2420 24980 2490
rect 24500 2370 24980 2420
rect 25640 1980 25880 3980
rect 7150 1740 25880 1980
rect -330 -140 150 -100
rect -330 -210 -300 -140
rect -230 -210 -190 -140
rect -120 -210 -80 -140
rect -10 -210 30 -140
rect 100 -210 150 -140
rect -330 -270 150 -210
rect -330 -340 -300 -270
rect -230 -340 -190 -270
rect -120 -340 -80 -270
rect -10 -340 30 -270
rect 100 -340 150 -270
rect -330 -380 150 -340
rect 7150 -120 7630 1740
rect 14590 1160 14900 1180
rect 14590 1090 14600 1160
rect 14670 1090 14700 1160
rect 14770 1090 14810 1160
rect 14880 1090 14900 1160
rect 14590 1050 14900 1090
rect 14590 980 14600 1050
rect 14670 980 14700 1050
rect 14770 980 14810 1050
rect 14880 980 14900 1050
rect 14590 940 14900 980
rect 14590 870 14600 940
rect 14670 870 14700 940
rect 14770 870 14810 940
rect 14880 870 14900 940
rect 14590 850 14900 870
rect 21060 920 21540 970
rect 21060 850 21090 920
rect 21160 850 21200 920
rect 21270 850 21310 920
rect 21380 850 21420 920
rect 21490 850 21540 920
rect 21060 810 21540 850
rect 21060 740 21090 810
rect 21160 740 21200 810
rect 21270 740 21310 810
rect 21380 740 21420 810
rect 21490 740 21540 810
rect 21060 710 21540 740
rect 23460 920 23940 970
rect 23460 850 23490 920
rect 23560 850 23600 920
rect 23670 850 23710 920
rect 23780 850 23820 920
rect 23890 850 23940 920
rect 23460 810 23940 850
rect 23460 740 23490 810
rect 23560 740 23600 810
rect 23670 740 23710 810
rect 23780 740 23820 810
rect 23890 740 23940 810
rect 23460 710 23940 740
rect 17040 0 28540 20
rect 17040 -20 28340 0
rect 17040 -90 20380 -20
rect 20450 -90 20490 -20
rect 20560 -90 20600 -20
rect 20670 -90 20710 -20
rect 20780 -70 28340 -20
rect 28410 -70 28450 0
rect 28520 -70 28540 0
rect 20780 -90 28540 -70
rect 7150 -180 7180 -120
rect 7240 -180 7280 -120
rect 7340 -180 7440 -120
rect 7500 -180 7540 -120
rect 7600 -180 7630 -120
rect 7150 -210 7630 -180
rect 7150 -270 7180 -210
rect 7240 -270 7280 -210
rect 7340 -270 7440 -210
rect 7500 -270 7540 -210
rect 7600 -270 7630 -210
rect 7150 -300 7630 -270
rect 7150 -360 7180 -300
rect 7240 -360 7280 -300
rect 7340 -360 7440 -300
rect 7500 -360 7540 -300
rect 7600 -360 7630 -300
rect 7150 -380 7630 -360
rect 14630 -140 15110 -100
rect 14630 -210 14660 -140
rect 14730 -210 14770 -140
rect 14840 -210 14880 -140
rect 14950 -210 14990 -140
rect 15060 -210 15110 -140
rect 14630 -270 15110 -210
rect 14630 -340 14660 -270
rect 14730 -340 14770 -270
rect 14840 -340 14880 -270
rect 14950 -340 14990 -270
rect 15060 -340 15110 -270
rect 14630 -380 15110 -340
rect 17040 -130 28540 -90
rect 17040 -200 20380 -130
rect 20450 -200 20490 -130
rect 20560 -200 20600 -130
rect 20670 -200 20710 -130
rect 20780 -200 28340 -130
rect 28410 -200 28450 -130
rect 28520 -200 28540 -130
rect 17040 -240 28540 -200
rect 17040 -310 20380 -240
rect 20450 -310 20490 -240
rect 20560 -310 20600 -240
rect 20670 -310 20710 -240
rect 20780 -260 28540 -240
rect 20780 -310 28340 -260
rect 17040 -330 28340 -310
rect 28410 -330 28450 -260
rect 28520 -330 28540 -260
rect 17040 -350 28540 -330
rect 1080 -790 2680 -760
rect 1080 -860 1150 -790
rect 1220 -860 1260 -790
rect 1330 -860 1370 -790
rect 1440 -860 1480 -790
rect 1550 -860 1590 -790
rect 1660 -860 1700 -790
rect 1770 -860 1810 -790
rect 1880 -860 1920 -790
rect 1990 -860 2030 -790
rect 2100 -860 2140 -790
rect 2210 -860 2250 -790
rect 2320 -860 2360 -790
rect 2430 -860 2470 -790
rect 2540 -860 2580 -790
rect 2650 -860 2680 -790
rect 1080 -900 2680 -860
rect 1080 -970 1150 -900
rect 1220 -970 1260 -900
rect 1330 -970 1370 -900
rect 1440 -970 1480 -900
rect 1550 -970 1590 -900
rect 1660 -970 1700 -900
rect 1770 -970 1810 -900
rect 1880 -970 1920 -900
rect 1990 -970 2030 -900
rect 2100 -970 2140 -900
rect 2210 -970 2250 -900
rect 2320 -970 2360 -900
rect 2430 -970 2470 -900
rect 2540 -970 2580 -900
rect 2650 -970 2680 -900
rect 1080 -1020 2680 -970
rect 12220 -790 13820 -760
rect 12220 -860 12250 -790
rect 12320 -860 12360 -790
rect 12430 -860 12470 -790
rect 12540 -860 12580 -790
rect 12650 -860 12690 -790
rect 12760 -860 12800 -790
rect 12870 -860 12910 -790
rect 12980 -860 13020 -790
rect 13090 -860 13130 -790
rect 13200 -860 13240 -790
rect 13310 -860 13350 -790
rect 13420 -860 13460 -790
rect 13530 -860 13570 -790
rect 13640 -860 13680 -790
rect 13750 -860 13820 -790
rect 12220 -900 13820 -860
rect 12220 -970 12250 -900
rect 12320 -970 12360 -900
rect 12430 -970 12470 -900
rect 12540 -970 12580 -900
rect 12650 -970 12690 -900
rect 12760 -970 12800 -900
rect 12870 -970 12910 -900
rect 12980 -970 13020 -900
rect 13090 -970 13130 -900
rect 13200 -970 13240 -900
rect 13310 -970 13350 -900
rect 13420 -970 13460 -900
rect 13530 -970 13570 -900
rect 13640 -970 13680 -900
rect 13750 -970 13820 -900
rect 12220 -1020 13820 -970
rect 1540 -2780 3140 -2730
rect 1540 -2850 1570 -2780
rect 1640 -2850 1680 -2780
rect 1750 -2850 1790 -2780
rect 1860 -2850 1900 -2780
rect 1970 -2850 2010 -2780
rect 2080 -2850 2120 -2780
rect 2190 -2850 2230 -2780
rect 2300 -2850 2340 -2780
rect 2410 -2850 2450 -2780
rect 2520 -2850 2560 -2780
rect 2630 -2850 2670 -2780
rect 2740 -2850 2780 -2780
rect 2850 -2850 2890 -2780
rect 2960 -2850 3000 -2780
rect 3070 -2850 3140 -2780
rect 1540 -2890 3140 -2850
rect 1540 -2960 1570 -2890
rect 1640 -2960 1680 -2890
rect 1750 -2960 1790 -2890
rect 1860 -2960 1900 -2890
rect 1970 -2960 2010 -2890
rect 2080 -2960 2120 -2890
rect 2190 -2960 2230 -2890
rect 2300 -2960 2340 -2890
rect 2410 -2960 2450 -2890
rect 2520 -2960 2560 -2890
rect 2630 -2960 2670 -2890
rect 2740 -2960 2780 -2890
rect 2850 -2960 2890 -2890
rect 2960 -2960 3000 -2890
rect 3070 -2960 3140 -2890
rect 1540 -2990 3140 -2960
rect 11760 -2780 13360 -2730
rect 11760 -2850 11790 -2780
rect 11860 -2850 11900 -2780
rect 11970 -2850 12010 -2780
rect 12080 -2850 12120 -2780
rect 12190 -2850 12230 -2780
rect 12300 -2850 12340 -2780
rect 12410 -2850 12450 -2780
rect 12520 -2850 12560 -2780
rect 12630 -2850 12670 -2780
rect 12740 -2850 12780 -2780
rect 12850 -2850 12890 -2780
rect 12960 -2850 13000 -2780
rect 13070 -2850 13110 -2780
rect 13180 -2850 13220 -2780
rect 13290 -2850 13360 -2780
rect 11760 -2890 13360 -2850
rect 11760 -2960 11790 -2890
rect 11860 -2960 11900 -2890
rect 11970 -2960 12010 -2890
rect 12080 -2960 12120 -2890
rect 12190 -2960 12230 -2890
rect 12300 -2960 12340 -2890
rect 12410 -2960 12450 -2890
rect 12520 -2960 12560 -2890
rect 12630 -2960 12670 -2890
rect 12740 -2960 12780 -2890
rect 12850 -2960 12890 -2890
rect 12960 -2960 13000 -2890
rect 13070 -2960 13110 -2890
rect 13180 -2960 13220 -2890
rect 13290 -2960 13360 -2890
rect 11760 -2990 13360 -2960
rect 17040 -3310 17280 -350
rect 25280 -1430 25880 -1400
rect 25280 -1490 25310 -1430
rect 25370 -1490 25410 -1430
rect 25470 -1490 25510 -1430
rect 25570 -1490 25880 -1430
rect 25280 -1530 25880 -1490
rect 25280 -1590 25310 -1530
rect 25370 -1590 25410 -1530
rect 25470 -1590 25510 -1530
rect 25570 -1590 25880 -1530
rect 25280 -1630 25880 -1590
rect 25280 -1690 25310 -1630
rect 25370 -1690 25410 -1630
rect 25470 -1690 25510 -1630
rect 25570 -1690 25880 -1630
rect 25280 -1730 25880 -1690
rect 25280 -1790 25310 -1730
rect 25370 -1790 25410 -1730
rect 25470 -1790 25510 -1730
rect 25570 -1790 25880 -1730
rect 25280 -1830 25880 -1790
rect 25280 -1890 25310 -1830
rect 25370 -1890 25410 -1830
rect 25470 -1890 25510 -1830
rect 25570 -1890 25880 -1830
rect 25280 -1930 25880 -1890
rect 25280 -1990 25310 -1930
rect 25370 -1990 25410 -1930
rect 25470 -1990 25510 -1930
rect 25570 -1990 25880 -1930
rect 25280 -2030 25880 -1990
rect 25280 -2090 25310 -2030
rect 25370 -2090 25410 -2030
rect 25470 -2090 25510 -2030
rect 25570 -2090 25880 -2030
rect 25280 -2130 25880 -2090
rect 25280 -2190 25310 -2130
rect 25370 -2190 25410 -2130
rect 25470 -2190 25510 -2130
rect 25570 -2190 25880 -2130
rect 25280 -2230 25880 -2190
rect 25280 -2290 25310 -2230
rect 25370 -2290 25410 -2230
rect 25470 -2290 25510 -2230
rect 25570 -2290 25880 -2230
rect 25280 -2320 25880 -2290
rect 7350 -3340 17280 -3310
rect 7350 -3400 7380 -3340
rect 7440 -3400 7480 -3340
rect 7540 -3400 17280 -3340
rect 22320 -3050 22650 -3030
rect 22320 -3120 22340 -3050
rect 22410 -3120 22450 -3050
rect 22520 -3120 22560 -3050
rect 22630 -3120 22650 -3050
rect 22320 -3160 22650 -3120
rect 22320 -3230 22340 -3160
rect 22410 -3230 22450 -3160
rect 22520 -3230 22560 -3160
rect 22630 -3230 22650 -3160
rect 22320 -3270 22650 -3230
rect 22320 -3340 22340 -3270
rect 22410 -3340 22450 -3270
rect 22520 -3340 22560 -3270
rect 22630 -3340 22650 -3270
rect 22320 -3360 22650 -3340
rect 7350 -3440 17280 -3400
rect 7350 -3550 7380 -3440
rect 7440 -3550 7480 -3440
rect 7540 -3550 17280 -3440
rect 7350 -3590 17280 -3550
rect 7350 -3650 7380 -3590
rect 7440 -3650 7480 -3590
rect 7540 -3650 17280 -3590
rect 7350 -3680 17280 -3650
rect 20020 -3690 20500 -3660
rect 20020 -3760 20070 -3690
rect 20140 -3760 20180 -3690
rect 20250 -3760 20290 -3690
rect 20360 -3760 20400 -3690
rect 20470 -3760 20500 -3690
rect 20020 -3800 20500 -3760
rect 20020 -3870 20070 -3800
rect 20140 -3870 20180 -3800
rect 20250 -3870 20290 -3800
rect 20360 -3870 20400 -3800
rect 20470 -3870 20500 -3800
rect 20020 -3920 20500 -3870
rect 24500 -3690 24980 -3660
rect 24500 -3760 24550 -3690
rect 24620 -3760 24660 -3690
rect 24730 -3760 24770 -3690
rect 24840 -3760 24880 -3690
rect 24950 -3760 24980 -3690
rect 24500 -3800 24980 -3760
rect 24500 -3870 24550 -3800
rect 24620 -3870 24660 -3800
rect 24730 -3870 24770 -3800
rect 24840 -3870 24880 -3800
rect 24950 -3870 24980 -3800
rect 24500 -3920 24980 -3870
rect 25680 -4370 25880 -2320
rect -2220 -4470 -2000 -4450
rect -2220 -4540 -2200 -4470
rect -2130 -4540 -2090 -4470
rect -2020 -4540 -2000 -4470
rect -2220 -4580 -2000 -4540
rect -2220 -4650 -2200 -4580
rect -2130 -4650 -2090 -4580
rect -2020 -4650 -2000 -4580
rect -2220 -4690 -2000 -4650
rect -2220 -4760 -2200 -4690
rect -2130 -4760 -2090 -4690
rect -2020 -4760 -2000 -4690
rect -2220 -4800 -2000 -4760
rect -2220 -4870 -2200 -4800
rect -2130 -4870 -2090 -4800
rect -2020 -4870 -2000 -4800
rect 7290 -4560 7620 -4540
rect 7290 -4630 7310 -4560
rect 7380 -4630 7420 -4560
rect 7490 -4630 7530 -4560
rect 7600 -4630 7620 -4560
rect 7290 -4670 7620 -4630
rect 7290 -4740 7310 -4670
rect 7380 -4740 7420 -4670
rect 7490 -4740 7530 -4670
rect 7600 -4740 7620 -4670
rect 7290 -4780 7620 -4740
rect 7290 -4850 7310 -4780
rect 7380 -4850 7420 -4780
rect 7490 -4850 7530 -4780
rect 7600 -4850 7620 -4780
rect 7290 -4870 7620 -4850
rect 17780 -4600 25880 -4370
rect -2220 -4890 -2000 -4870
rect -2160 -5240 -1940 -5220
rect -2160 -5310 -2140 -5240
rect -2070 -5310 -2030 -5240
rect -1960 -5310 -1940 -5240
rect -2160 -5350 -1940 -5310
rect -2160 -5420 -2140 -5350
rect -2070 -5420 -2030 -5350
rect -1960 -5420 -1940 -5350
rect -2160 -5460 -1940 -5420
rect -2160 -5530 -2140 -5460
rect -2070 -5530 -2030 -5460
rect -1960 -5530 -1940 -5460
rect -2160 -5570 -1940 -5530
rect -2160 -5640 -2140 -5570
rect -2070 -5640 -2030 -5570
rect -1960 -5640 -1940 -5570
rect -2160 -5660 -1940 -5640
rect 7030 -6460 7340 -6420
rect -880 -6500 -600 -6470
rect -880 -6570 -840 -6500
rect -770 -6570 -710 -6500
rect -640 -6570 -600 -6500
rect -880 -6610 -600 -6570
rect -880 -6680 -840 -6610
rect -770 -6680 -710 -6610
rect -640 -6680 -600 -6610
rect 7030 -6520 7050 -6460
rect 7110 -6520 7150 -6460
rect 7210 -6520 7250 -6460
rect 7310 -6520 7340 -6460
rect 7030 -6560 7340 -6520
rect 7030 -6620 7050 -6560
rect 7110 -6620 7150 -6560
rect 7210 -6620 7250 -6560
rect 7310 -6620 7340 -6560
rect -880 -6720 -600 -6680
rect -880 -6790 -840 -6720
rect -770 -6790 -710 -6720
rect -640 -6790 -600 -6720
rect -880 -6830 -600 -6790
rect -880 -6900 -840 -6830
rect -770 -6900 -710 -6830
rect -640 -6900 -600 -6830
rect -880 -6950 -600 -6900
rect 4740 -6670 5060 -6640
rect 4740 -6730 4770 -6670
rect 4830 -6730 4870 -6670
rect 4930 -6730 4970 -6670
rect 5030 -6730 5060 -6670
rect 4740 -6770 5060 -6730
rect 4740 -6830 4770 -6770
rect 4830 -6830 4870 -6770
rect 4930 -6830 4970 -6770
rect 5030 -6830 5060 -6770
rect 4740 -6870 5060 -6830
rect 7030 -6660 7340 -6620
rect 7030 -6720 7050 -6660
rect 7110 -6720 7150 -6660
rect 7210 -6720 7250 -6660
rect 7310 -6720 7340 -6660
rect 7030 -6760 7340 -6720
rect 7030 -6820 7050 -6760
rect 7110 -6820 7150 -6760
rect 7210 -6820 7250 -6760
rect 7310 -6820 7340 -6760
rect 7030 -6850 7340 -6820
rect 7570 -6460 7870 -6420
rect 7570 -6520 7590 -6460
rect 7650 -6520 7690 -6460
rect 7750 -6520 7790 -6460
rect 7850 -6520 7870 -6460
rect 7570 -6560 7870 -6520
rect 7570 -6620 7590 -6560
rect 7650 -6620 7690 -6560
rect 7750 -6620 7790 -6560
rect 7850 -6620 7870 -6560
rect 7570 -6660 7870 -6620
rect 15380 -6500 15660 -6470
rect 15380 -6570 15420 -6500
rect 15490 -6570 15550 -6500
rect 15620 -6570 15660 -6500
rect 15380 -6610 15660 -6570
rect 7570 -6720 7590 -6660
rect 7650 -6720 7690 -6660
rect 7750 -6720 7790 -6660
rect 7850 -6720 7870 -6660
rect 7570 -6760 7870 -6720
rect 7570 -6820 7590 -6760
rect 7650 -6820 7690 -6760
rect 7750 -6820 7790 -6760
rect 7850 -6820 7870 -6760
rect 7570 -6850 7870 -6820
rect 9840 -6670 10160 -6640
rect 9840 -6730 9870 -6670
rect 9930 -6730 9970 -6670
rect 10030 -6730 10070 -6670
rect 10130 -6730 10160 -6670
rect 9840 -6770 10160 -6730
rect 9840 -6830 9870 -6770
rect 9930 -6830 9970 -6770
rect 10030 -6830 10070 -6770
rect 10130 -6830 10160 -6770
rect 4740 -6930 4770 -6870
rect 4830 -6930 4870 -6870
rect 4930 -6930 4970 -6870
rect 5030 -6930 5060 -6870
rect 4740 -6950 5060 -6930
rect 9840 -6870 10160 -6830
rect 9840 -6930 9870 -6870
rect 9930 -6930 9970 -6870
rect 10030 -6930 10070 -6870
rect 10130 -6930 10160 -6870
rect 9840 -6950 10160 -6930
rect 15380 -6680 15420 -6610
rect 15490 -6680 15550 -6610
rect 15620 -6680 15660 -6610
rect 15380 -6720 15660 -6680
rect 15380 -6790 15420 -6720
rect 15490 -6790 15550 -6720
rect 15620 -6790 15660 -6720
rect 15380 -6830 15660 -6790
rect 15380 -6900 15420 -6830
rect 15490 -6900 15550 -6830
rect 15620 -6900 15660 -6830
rect 15380 -6950 15660 -6900
rect -2220 -7870 -2000 -7850
rect -2220 -7940 -2200 -7870
rect -2130 -7940 -2090 -7870
rect -2020 -7940 -2000 -7870
rect -2220 -7980 -2000 -7940
rect -2220 -8050 -2200 -7980
rect -2130 -8050 -2090 -7980
rect -2020 -8050 -2000 -7980
rect -2220 -8090 -2000 -8050
rect -2220 -8160 -2200 -8090
rect -2130 -8160 -2090 -8090
rect -2020 -8160 -2000 -8090
rect -2220 -8200 -2000 -8160
rect -2220 -8270 -2200 -8200
rect -2130 -8270 -2090 -8200
rect -2020 -8270 -2000 -8200
rect -2220 -8290 -2000 -8270
rect 14590 -8230 14900 -8210
rect 14590 -8300 14600 -8230
rect 14670 -8300 14700 -8230
rect 14770 -8300 14810 -8230
rect 14880 -8300 14900 -8230
rect 14590 -8340 14900 -8300
rect 14590 -8410 14600 -8340
rect 14670 -8410 14700 -8340
rect 14770 -8410 14810 -8340
rect 14880 -8410 14900 -8340
rect 14590 -8450 14900 -8410
rect 14590 -8520 14600 -8450
rect 14670 -8520 14700 -8450
rect 14770 -8520 14810 -8450
rect 14880 -8520 14900 -8450
rect 14590 -8540 14900 -8520
rect -2160 -8640 -1940 -8620
rect -2160 -8710 -2140 -8640
rect -2070 -8710 -2030 -8640
rect -1960 -8710 -1940 -8640
rect -2160 -8750 -1940 -8710
rect -2160 -8820 -2140 -8750
rect -2070 -8820 -2030 -8750
rect -1960 -8820 -1940 -8750
rect -2160 -8860 -1940 -8820
rect -2160 -8930 -2140 -8860
rect -2070 -8930 -2030 -8860
rect -1960 -8930 -1940 -8860
rect -2160 -8970 -1940 -8930
rect -2160 -9040 -2140 -8970
rect -2070 -9040 -2030 -8970
rect -1960 -9040 -1940 -8970
rect -2160 -9060 -1940 -9040
rect 17780 -9160 18090 -4600
rect 19210 -8560 19530 -8530
rect 19210 -8630 19230 -8560
rect 19300 -8630 19330 -8560
rect 19400 -8630 19430 -8560
rect 19500 -8630 19530 -8560
rect 19210 -8660 19530 -8630
rect 19210 -8730 19230 -8660
rect 19300 -8730 19330 -8660
rect 19400 -8730 19430 -8660
rect 19500 -8730 19530 -8660
rect 19210 -8760 19530 -8730
rect 19210 -8830 19230 -8760
rect 19300 -8830 19330 -8760
rect 19400 -8830 19430 -8760
rect 19500 -8830 19530 -8760
rect 19210 -8850 19530 -8830
rect 7210 -9440 18090 -9160
rect 19940 -9000 20260 -8970
rect 19940 -9070 19960 -9000
rect 20030 -9070 20060 -9000
rect 20130 -9070 20160 -9000
rect 20230 -9070 20260 -9000
rect 19940 -9100 20260 -9070
rect 19940 -9170 19960 -9100
rect 20030 -9170 20060 -9100
rect 20130 -9170 20160 -9100
rect 20230 -9170 20260 -9100
rect 19940 -9200 20260 -9170
rect 19940 -9270 19960 -9200
rect 20030 -9270 20060 -9200
rect 20130 -9270 20160 -9200
rect 20230 -9270 20260 -9200
rect 19940 -9290 20260 -9270
rect -270 -9660 210 -9620
rect -270 -9730 -240 -9660
rect -170 -9730 -130 -9660
rect -60 -9730 -20 -9660
rect 50 -9730 90 -9660
rect 160 -9730 210 -9660
rect -270 -9790 210 -9730
rect -270 -9860 -240 -9790
rect -170 -9860 -130 -9790
rect -60 -9860 -20 -9790
rect 50 -9860 90 -9790
rect 160 -9860 210 -9790
rect -270 -9900 210 -9860
rect 7210 -9640 7690 -9440
rect 7210 -9700 7240 -9640
rect 7300 -9700 7340 -9640
rect 7400 -9700 7500 -9640
rect 7560 -9700 7600 -9640
rect 7660 -9700 7690 -9640
rect 7210 -9730 7690 -9700
rect 7210 -9790 7240 -9730
rect 7300 -9790 7340 -9730
rect 7400 -9790 7500 -9730
rect 7560 -9790 7600 -9730
rect 7660 -9790 7690 -9730
rect 7210 -9820 7690 -9790
rect 7210 -9880 7240 -9820
rect 7300 -9880 7340 -9820
rect 7400 -9880 7500 -9820
rect 7560 -9880 7600 -9820
rect 7660 -9880 7690 -9820
rect 7210 -9900 7690 -9880
rect 14690 -9660 15170 -9620
rect 14690 -9730 14720 -9660
rect 14790 -9730 14830 -9660
rect 14900 -9730 14940 -9660
rect 15010 -9730 15050 -9660
rect 15120 -9730 15170 -9660
rect 14690 -9790 15170 -9730
rect 14690 -9860 14720 -9790
rect 14790 -9860 14830 -9790
rect 14900 -9860 14940 -9790
rect 15010 -9860 15050 -9790
rect 15120 -9860 15170 -9790
rect 14690 -9900 15170 -9860
rect 1080 -10340 2680 -10310
rect 1080 -10410 1150 -10340
rect 1220 -10410 1260 -10340
rect 1330 -10410 1370 -10340
rect 1440 -10410 1480 -10340
rect 1550 -10410 1590 -10340
rect 1660 -10410 1700 -10340
rect 1770 -10410 1810 -10340
rect 1880 -10410 1920 -10340
rect 1990 -10410 2030 -10340
rect 2100 -10410 2140 -10340
rect 2210 -10410 2250 -10340
rect 2320 -10410 2360 -10340
rect 2430 -10410 2470 -10340
rect 2540 -10410 2580 -10340
rect 2650 -10410 2680 -10340
rect 1080 -10450 2680 -10410
rect 1080 -10520 1150 -10450
rect 1220 -10520 1260 -10450
rect 1330 -10520 1370 -10450
rect 1440 -10520 1480 -10450
rect 1550 -10520 1590 -10450
rect 1660 -10520 1700 -10450
rect 1770 -10520 1810 -10450
rect 1880 -10520 1920 -10450
rect 1990 -10520 2030 -10450
rect 2100 -10520 2140 -10450
rect 2210 -10520 2250 -10450
rect 2320 -10520 2360 -10450
rect 2430 -10520 2470 -10450
rect 2540 -10520 2580 -10450
rect 2650 -10520 2680 -10450
rect 1080 -10570 2680 -10520
rect 12220 -10370 13820 -10340
rect 12220 -10440 12290 -10370
rect 12360 -10440 12400 -10370
rect 12470 -10440 12510 -10370
rect 12580 -10440 12620 -10370
rect 12690 -10440 12730 -10370
rect 12800 -10440 12840 -10370
rect 12910 -10440 12950 -10370
rect 13020 -10440 13060 -10370
rect 13130 -10440 13170 -10370
rect 13240 -10440 13280 -10370
rect 13350 -10440 13390 -10370
rect 13460 -10440 13500 -10370
rect 13570 -10440 13610 -10370
rect 13680 -10440 13720 -10370
rect 13790 -10440 13820 -10370
rect 12220 -10480 13820 -10440
rect 12220 -10550 12290 -10480
rect 12360 -10550 12400 -10480
rect 12470 -10550 12510 -10480
rect 12580 -10550 12620 -10480
rect 12690 -10550 12730 -10480
rect 12800 -10550 12840 -10480
rect 12910 -10550 12950 -10480
rect 13020 -10550 13060 -10480
rect 13130 -10550 13170 -10480
rect 13240 -10550 13280 -10480
rect 13350 -10550 13390 -10480
rect 13460 -10550 13500 -10480
rect 13570 -10550 13610 -10480
rect 13680 -10550 13720 -10480
rect 13790 -10550 13820 -10480
rect 12220 -10600 13820 -10550
rect 2210 -12300 3810 -12250
rect 2210 -12370 2240 -12300
rect 2310 -12370 2350 -12300
rect 2420 -12370 2460 -12300
rect 2530 -12370 2570 -12300
rect 2640 -12370 2680 -12300
rect 2750 -12370 2790 -12300
rect 2860 -12370 2900 -12300
rect 2970 -12370 3010 -12300
rect 3080 -12370 3120 -12300
rect 3190 -12370 3230 -12300
rect 3300 -12370 3340 -12300
rect 3410 -12370 3450 -12300
rect 3520 -12370 3560 -12300
rect 3630 -12370 3670 -12300
rect 3740 -12370 3810 -12300
rect 2210 -12410 3810 -12370
rect 2210 -12480 2240 -12410
rect 2310 -12480 2350 -12410
rect 2420 -12480 2460 -12410
rect 2530 -12480 2570 -12410
rect 2640 -12480 2680 -12410
rect 2750 -12480 2790 -12410
rect 2860 -12480 2900 -12410
rect 2970 -12480 3010 -12410
rect 3080 -12480 3120 -12410
rect 3190 -12480 3230 -12410
rect 3300 -12480 3340 -12410
rect 3410 -12480 3450 -12410
rect 3520 -12480 3560 -12410
rect 3630 -12480 3670 -12410
rect 3740 -12480 3810 -12410
rect 2210 -12510 3810 -12480
rect 11090 -12300 12690 -12250
rect 11090 -12370 11120 -12300
rect 11190 -12370 11230 -12300
rect 11300 -12370 11340 -12300
rect 11410 -12370 11450 -12300
rect 11520 -12370 11560 -12300
rect 11630 -12370 11670 -12300
rect 11740 -12370 11780 -12300
rect 11850 -12370 11890 -12300
rect 11960 -12370 12000 -12300
rect 12070 -12370 12110 -12300
rect 12180 -12370 12220 -12300
rect 12290 -12370 12330 -12300
rect 12400 -12370 12440 -12300
rect 12510 -12370 12550 -12300
rect 12620 -12370 12690 -12300
rect 11090 -12410 12690 -12370
rect 11090 -12480 11120 -12410
rect 11190 -12480 11230 -12410
rect 11300 -12480 11340 -12410
rect 11410 -12480 11450 -12410
rect 11520 -12480 11560 -12410
rect 11630 -12480 11670 -12410
rect 11740 -12480 11780 -12410
rect 11850 -12480 11890 -12410
rect 11960 -12480 12000 -12410
rect 12070 -12480 12110 -12410
rect 12180 -12480 12220 -12410
rect 12290 -12480 12330 -12410
rect 12400 -12480 12440 -12410
rect 12510 -12480 12550 -12410
rect 12620 -12480 12690 -12410
rect 11090 -12510 12690 -12480
rect 6980 -13250 7310 -13220
rect 6980 -13310 7010 -13250
rect 7070 -13310 7110 -13250
rect 7170 -13310 7210 -13250
rect 7270 -13310 7310 -13250
rect 6980 -13340 7310 -13310
rect 6980 -13400 7010 -13340
rect 7070 -13400 7110 -13340
rect 7170 -13400 7210 -13340
rect 7270 -13400 7310 -13340
rect 6980 -13430 7310 -13400
rect 6980 -13490 7010 -13430
rect 7070 -13490 7110 -13430
rect 7170 -13490 7210 -13430
rect 7270 -13490 7310 -13430
rect 6980 -13530 7310 -13490
rect 6980 -13590 7010 -13530
rect 7070 -13590 7110 -13530
rect 7170 -13590 7210 -13530
rect 7270 -13590 7310 -13530
rect 6980 -13620 7310 -13590
rect 6980 -13680 7010 -13620
rect 7070 -13680 7110 -13620
rect 7170 -13680 7210 -13620
rect 7270 -13680 7310 -13620
rect 6980 -13710 7310 -13680
rect 6980 -13770 7010 -13710
rect 7070 -13770 7110 -13710
rect 7170 -13770 7210 -13710
rect 7270 -13770 7310 -13710
rect 6980 -13800 7310 -13770
rect 7590 -13250 7920 -13220
rect 7590 -13310 7630 -13250
rect 7690 -13310 7730 -13250
rect 7790 -13310 7830 -13250
rect 7890 -13310 7920 -13250
rect 7590 -13340 7920 -13310
rect 7590 -13400 7630 -13340
rect 7690 -13400 7730 -13340
rect 7790 -13400 7830 -13340
rect 7890 -13400 7920 -13340
rect 7590 -13430 7920 -13400
rect 7590 -13490 7630 -13430
rect 7690 -13490 7730 -13430
rect 7790 -13490 7830 -13430
rect 7890 -13490 7920 -13430
rect 7590 -13530 7920 -13490
rect 7590 -13590 7630 -13530
rect 7690 -13590 7730 -13530
rect 7790 -13590 7830 -13530
rect 7890 -13590 7920 -13530
rect 7590 -13620 7920 -13590
rect 7590 -13680 7630 -13620
rect 7690 -13680 7730 -13620
rect 7790 -13680 7830 -13620
rect 7890 -13680 7920 -13620
rect 7590 -13710 7920 -13680
rect 7590 -13770 7630 -13710
rect 7690 -13770 7730 -13710
rect 7790 -13770 7830 -13710
rect 7890 -13770 7920 -13710
rect 7590 -13800 7920 -13770
rect 19210 -14220 19530 -14190
rect 19210 -14290 19230 -14220
rect 19300 -14290 19330 -14220
rect 19400 -14290 19430 -14220
rect 19500 -14290 19530 -14220
rect 19210 -14320 19530 -14290
rect 19210 -14390 19230 -14320
rect 19300 -14390 19330 -14320
rect 19400 -14390 19430 -14320
rect 19500 -14390 19530 -14320
rect 19210 -14420 19530 -14390
rect 19210 -14490 19230 -14420
rect 19300 -14490 19330 -14420
rect 19400 -14490 19430 -14420
rect 19500 -14490 19530 -14420
rect 19210 -14510 19530 -14490
rect 20460 -14870 20780 -14840
rect 20460 -14940 20480 -14870
rect 20550 -14940 20580 -14870
rect 20650 -14940 20680 -14870
rect 20750 -14940 20780 -14870
rect 20460 -14970 20780 -14940
rect 20460 -15040 20480 -14970
rect 20550 -15040 20580 -14970
rect 20650 -15040 20680 -14970
rect 20750 -15040 20780 -14970
rect 20460 -15070 20780 -15040
rect 20460 -15140 20480 -15070
rect 20550 -15140 20580 -15070
rect 20650 -15140 20680 -15070
rect 20750 -15140 20780 -15070
rect 20460 -15160 20780 -15140
rect 5010 -17100 5330 -17070
rect 5010 -17160 5040 -17100
rect 5100 -17160 5140 -17100
rect 5200 -17160 5240 -17100
rect 5300 -17160 5330 -17100
rect 5010 -17200 5330 -17160
rect 5010 -17260 5040 -17200
rect 5100 -17260 5140 -17200
rect 5200 -17260 5240 -17200
rect 5300 -17260 5330 -17200
rect 5010 -17300 5330 -17260
rect 5010 -17360 5040 -17300
rect 5100 -17360 5140 -17300
rect 5200 -17360 5240 -17300
rect 5300 -17360 5330 -17300
rect 5010 -17380 5330 -17360
rect 9570 -17100 9890 -17070
rect 9570 -17160 9600 -17100
rect 9660 -17160 9700 -17100
rect 9760 -17160 9800 -17100
rect 9860 -17160 9890 -17100
rect 9570 -17200 9890 -17160
rect 9570 -17260 9600 -17200
rect 9660 -17260 9700 -17200
rect 9760 -17260 9800 -17200
rect 9860 -17260 9890 -17200
rect 9570 -17300 9890 -17260
rect 9570 -17360 9600 -17300
rect 9660 -17360 9700 -17300
rect 9760 -17360 9800 -17300
rect 9860 -17360 9890 -17300
rect 9570 -17380 9890 -17360
rect 7210 -17600 7650 -17580
rect 7210 -17670 7230 -17600
rect 7300 -17670 7340 -17600
rect 7410 -17670 7450 -17600
rect 7520 -17670 7560 -17600
rect 7630 -17670 7650 -17600
rect 7210 -17710 7650 -17670
rect 7210 -17780 7230 -17710
rect 7300 -17780 7340 -17710
rect 7410 -17780 7450 -17710
rect 7520 -17780 7560 -17710
rect 7630 -17780 7650 -17710
rect 7210 -17820 7650 -17780
rect 7210 -17890 7230 -17820
rect 7300 -17890 7340 -17820
rect 7410 -17890 7450 -17820
rect 7520 -17890 7560 -17820
rect 7630 -17890 7650 -17820
rect 7210 -17930 7650 -17890
rect 7210 -18000 7230 -17930
rect 7300 -18000 7340 -17930
rect 7410 -18000 7450 -17930
rect 7520 -18000 7560 -17930
rect 7630 -18000 7650 -17930
rect 7210 -18020 7650 -18000
rect 19210 -20290 19530 -20260
rect 19210 -20360 19230 -20290
rect 19300 -20360 19330 -20290
rect 19400 -20360 19430 -20290
rect 19500 -20360 19530 -20290
rect 19210 -20390 19530 -20360
rect 19210 -20460 19230 -20390
rect 19300 -20460 19330 -20390
rect 19400 -20460 19430 -20390
rect 19500 -20460 19530 -20390
rect 19210 -20490 19530 -20460
rect 19210 -20560 19230 -20490
rect 19300 -20560 19330 -20490
rect 19400 -20560 19430 -20490
rect 19500 -20560 19530 -20490
rect 19210 -20580 19530 -20560
rect 20020 -20720 20340 -20690
rect 20020 -20790 20040 -20720
rect 20110 -20790 20140 -20720
rect 20210 -20790 20240 -20720
rect 20310 -20790 20340 -20720
rect 20020 -20820 20340 -20790
rect 20020 -20890 20040 -20820
rect 20110 -20890 20140 -20820
rect 20210 -20890 20240 -20820
rect 20310 -20890 20340 -20820
rect 20020 -20920 20340 -20890
rect 20020 -20990 20040 -20920
rect 20110 -20990 20140 -20920
rect 20210 -20990 20240 -20920
rect 20310 -20990 20340 -20920
rect 20020 -21010 20340 -20990
rect 2210 -22660 3810 -22630
rect 2210 -22730 2280 -22660
rect 2350 -22730 2390 -22660
rect 2460 -22730 2500 -22660
rect 2570 -22730 2610 -22660
rect 2680 -22730 2720 -22660
rect 2790 -22730 2830 -22660
rect 2900 -22730 2940 -22660
rect 3010 -22730 3050 -22660
rect 3120 -22730 3160 -22660
rect 3230 -22730 3270 -22660
rect 3340 -22730 3380 -22660
rect 3450 -22730 3490 -22660
rect 3560 -22730 3600 -22660
rect 3670 -22730 3710 -22660
rect 3780 -22730 3810 -22660
rect 2210 -22770 3810 -22730
rect 2210 -22840 2280 -22770
rect 2350 -22840 2390 -22770
rect 2460 -22840 2500 -22770
rect 2570 -22840 2610 -22770
rect 2680 -22840 2720 -22770
rect 2790 -22840 2830 -22770
rect 2900 -22840 2940 -22770
rect 3010 -22840 3050 -22770
rect 3120 -22840 3160 -22770
rect 3230 -22840 3270 -22770
rect 3340 -22840 3380 -22770
rect 3450 -22840 3490 -22770
rect 3560 -22840 3600 -22770
rect 3670 -22840 3710 -22770
rect 3780 -22840 3810 -22770
rect 2210 -22890 3810 -22840
rect 11090 -22660 12690 -22630
rect 11090 -22730 11160 -22660
rect 11230 -22730 11270 -22660
rect 11340 -22730 11380 -22660
rect 11450 -22730 11490 -22660
rect 11560 -22730 11600 -22660
rect 11670 -22730 11710 -22660
rect 11780 -22730 11820 -22660
rect 11890 -22730 11930 -22660
rect 12000 -22730 12040 -22660
rect 12110 -22730 12150 -22660
rect 12220 -22730 12260 -22660
rect 12330 -22730 12370 -22660
rect 12440 -22730 12480 -22660
rect 12550 -22730 12590 -22660
rect 12660 -22730 12690 -22660
rect 11090 -22770 12690 -22730
rect 11090 -22840 11160 -22770
rect 11230 -22840 11270 -22770
rect 11340 -22840 11380 -22770
rect 11450 -22840 11490 -22770
rect 11560 -22840 11600 -22770
rect 11670 -22840 11710 -22770
rect 11780 -22840 11820 -22770
rect 11890 -22840 11930 -22770
rect 12000 -22840 12040 -22770
rect 12110 -22840 12150 -22770
rect 12220 -22840 12260 -22770
rect 12330 -22840 12370 -22770
rect 12440 -22840 12480 -22770
rect 12550 -22840 12590 -22770
rect 12660 -22840 12690 -22770
rect 11090 -22890 12690 -22840
<< via2 >>
rect 21090 7140 21160 7210
rect 21200 7140 21270 7210
rect 21310 7140 21380 7210
rect 21420 7140 21490 7210
rect 21090 7030 21160 7100
rect 21200 7030 21270 7100
rect 21310 7030 21380 7100
rect 21420 7030 21490 7100
rect 23490 7140 23560 7210
rect 23600 7140 23670 7210
rect 23710 7140 23780 7210
rect 23820 7140 23890 7210
rect 23490 7030 23560 7100
rect 23600 7030 23670 7100
rect 23710 7030 23780 7100
rect 23820 7030 23890 7100
rect 1570 6780 1640 6850
rect 1680 6780 1750 6850
rect 1790 6780 1860 6850
rect 1900 6780 1970 6850
rect 2010 6780 2080 6850
rect 2120 6780 2190 6850
rect 2230 6780 2300 6850
rect 2340 6780 2410 6850
rect 2450 6780 2520 6850
rect 2560 6780 2630 6850
rect 2670 6780 2740 6850
rect 2780 6780 2850 6850
rect 2890 6780 2960 6850
rect 3000 6780 3070 6850
rect 1570 6670 1640 6740
rect 1680 6670 1750 6740
rect 1790 6670 1860 6740
rect 1900 6670 1970 6740
rect 2010 6670 2080 6740
rect 2120 6670 2190 6740
rect 2230 6670 2300 6740
rect 2340 6670 2410 6740
rect 2450 6670 2520 6740
rect 2560 6670 2630 6740
rect 2670 6670 2740 6740
rect 2780 6670 2850 6740
rect 2890 6670 2960 6740
rect 3000 6670 3070 6740
rect 11790 6810 11860 6880
rect 11900 6810 11970 6880
rect 12010 6810 12080 6880
rect 12120 6810 12190 6880
rect 12230 6810 12300 6880
rect 12340 6810 12410 6880
rect 12450 6810 12520 6880
rect 12560 6810 12630 6880
rect 12670 6810 12740 6880
rect 12780 6810 12850 6880
rect 12890 6810 12960 6880
rect 13000 6810 13070 6880
rect 13110 6810 13180 6880
rect 13220 6810 13290 6880
rect 11790 6700 11860 6770
rect 11900 6700 11970 6770
rect 12010 6700 12080 6770
rect 12120 6700 12190 6770
rect 12230 6700 12300 6770
rect 12340 6700 12410 6770
rect 12450 6700 12520 6770
rect 12560 6700 12630 6770
rect 12670 6700 12740 6770
rect 12780 6700 12850 6770
rect 12890 6700 12960 6770
rect 13000 6700 13070 6770
rect 13110 6700 13180 6770
rect 13220 6700 13290 6770
rect 28340 6230 28410 6300
rect 28450 6230 28520 6300
rect 28340 6100 28410 6170
rect 28450 6100 28520 6170
rect 28340 5970 28410 6040
rect 28450 5970 28520 6040
rect 7410 5320 7480 5390
rect 7410 5210 7480 5280
rect 7410 5100 7480 5170
rect 7410 4990 7480 5060
rect 7410 4880 7480 4950
rect 7590 4700 7650 4760
rect 7690 4700 7750 4760
rect 7790 4700 7850 4760
rect -840 4510 -770 4580
rect -710 4510 -640 4580
rect -840 4400 -770 4470
rect -710 4400 -640 4470
rect -840 4290 -770 4360
rect -710 4290 -640 4360
rect -840 4180 -770 4250
rect -710 4180 -640 4250
rect 6700 4520 6760 4580
rect 6700 4400 6760 4460
rect 6700 4280 6760 4340
rect 6700 4160 6760 4220
rect 15420 4510 15490 4580
rect 15550 4510 15620 4580
rect 15420 4400 15490 4470
rect 15550 4400 15620 4470
rect 15420 4290 15490 4360
rect 15550 4290 15620 4360
rect 15420 4180 15490 4250
rect 15550 4180 15620 4250
rect 7050 3180 7110 3240
rect 7150 3180 7210 3240
rect 7250 3180 7310 3240
rect 7050 3080 7110 3140
rect 7150 3080 7210 3140
rect 7250 3080 7310 3140
rect 7050 2980 7110 3040
rect 7150 2980 7210 3040
rect 7250 2980 7310 3040
rect 22320 3290 22390 3360
rect 22430 3290 22500 3360
rect 22540 3290 22610 3360
rect 22320 3180 22390 3250
rect 22430 3180 22500 3250
rect 22540 3180 22610 3250
rect 22320 3070 22390 3140
rect 22430 3070 22500 3140
rect 22540 3070 22610 3140
rect 4770 2830 4830 2890
rect 4870 2830 4930 2890
rect 4970 2830 5030 2890
rect 4770 2730 4830 2790
rect 4870 2730 4930 2790
rect 4970 2730 5030 2790
rect 4770 2630 4830 2690
rect 4870 2630 4930 2690
rect 4970 2630 5030 2690
rect 9870 2830 9930 2890
rect 9970 2830 10030 2890
rect 10070 2830 10130 2890
rect 9870 2730 9930 2790
rect 9970 2730 10030 2790
rect 10070 2730 10130 2790
rect 9870 2630 9930 2690
rect 9970 2630 10030 2690
rect 10070 2630 10130 2690
rect 20070 2530 20140 2600
rect 20180 2530 20250 2600
rect 20290 2530 20360 2600
rect 20400 2530 20470 2600
rect 20070 2420 20140 2490
rect 20180 2420 20250 2490
rect 20290 2420 20360 2490
rect 20400 2420 20470 2490
rect 24550 2530 24620 2600
rect 24660 2530 24730 2600
rect 24770 2530 24840 2600
rect 24880 2530 24950 2600
rect 24550 2420 24620 2490
rect 24660 2420 24730 2490
rect 24770 2420 24840 2490
rect 24880 2420 24950 2490
rect -300 -210 -230 -140
rect -190 -210 -120 -140
rect -80 -210 -10 -140
rect 30 -210 100 -140
rect -300 -340 -230 -270
rect -190 -340 -120 -270
rect -80 -340 -10 -270
rect 30 -340 100 -270
rect 14600 1090 14670 1160
rect 14700 1090 14770 1160
rect 14810 1090 14880 1160
rect 14600 980 14670 1050
rect 14700 980 14770 1050
rect 14810 980 14880 1050
rect 14600 870 14670 940
rect 14700 870 14770 940
rect 14810 870 14880 940
rect 21090 850 21160 920
rect 21200 850 21270 920
rect 21310 850 21380 920
rect 21420 850 21490 920
rect 21090 740 21160 810
rect 21200 740 21270 810
rect 21310 740 21380 810
rect 21420 740 21490 810
rect 23490 850 23560 920
rect 23600 850 23670 920
rect 23710 850 23780 920
rect 23820 850 23890 920
rect 23490 740 23560 810
rect 23600 740 23670 810
rect 23710 740 23780 810
rect 23820 740 23890 810
rect 28340 -70 28410 0
rect 28450 -70 28520 0
rect 14660 -210 14730 -140
rect 14770 -210 14840 -140
rect 14880 -210 14950 -140
rect 14990 -210 15060 -140
rect 14660 -340 14730 -270
rect 14770 -340 14840 -270
rect 14880 -340 14950 -270
rect 14990 -340 15060 -270
rect 28340 -200 28410 -130
rect 28450 -200 28520 -130
rect 28340 -330 28410 -260
rect 28450 -330 28520 -260
rect 1150 -860 1220 -790
rect 1260 -860 1330 -790
rect 1370 -860 1440 -790
rect 1480 -860 1550 -790
rect 1590 -860 1660 -790
rect 1700 -860 1770 -790
rect 1810 -860 1880 -790
rect 1920 -860 1990 -790
rect 2030 -860 2100 -790
rect 2140 -860 2210 -790
rect 2250 -860 2320 -790
rect 2360 -860 2430 -790
rect 2470 -860 2540 -790
rect 2580 -860 2650 -790
rect 1150 -970 1220 -900
rect 1260 -970 1330 -900
rect 1370 -970 1440 -900
rect 1480 -970 1550 -900
rect 1590 -970 1660 -900
rect 1700 -970 1770 -900
rect 1810 -970 1880 -900
rect 1920 -970 1990 -900
rect 2030 -970 2100 -900
rect 2140 -970 2210 -900
rect 2250 -970 2320 -900
rect 2360 -970 2430 -900
rect 2470 -970 2540 -900
rect 2580 -970 2650 -900
rect 12250 -860 12320 -790
rect 12360 -860 12430 -790
rect 12470 -860 12540 -790
rect 12580 -860 12650 -790
rect 12690 -860 12760 -790
rect 12800 -860 12870 -790
rect 12910 -860 12980 -790
rect 13020 -860 13090 -790
rect 13130 -860 13200 -790
rect 13240 -860 13310 -790
rect 13350 -860 13420 -790
rect 13460 -860 13530 -790
rect 13570 -860 13640 -790
rect 13680 -860 13750 -790
rect 12250 -970 12320 -900
rect 12360 -970 12430 -900
rect 12470 -970 12540 -900
rect 12580 -970 12650 -900
rect 12690 -970 12760 -900
rect 12800 -970 12870 -900
rect 12910 -970 12980 -900
rect 13020 -970 13090 -900
rect 13130 -970 13200 -900
rect 13240 -970 13310 -900
rect 13350 -970 13420 -900
rect 13460 -970 13530 -900
rect 13570 -970 13640 -900
rect 13680 -970 13750 -900
rect 1570 -2850 1640 -2780
rect 1680 -2850 1750 -2780
rect 1790 -2850 1860 -2780
rect 1900 -2850 1970 -2780
rect 2010 -2850 2080 -2780
rect 2120 -2850 2190 -2780
rect 2230 -2850 2300 -2780
rect 2340 -2850 2410 -2780
rect 2450 -2850 2520 -2780
rect 2560 -2850 2630 -2780
rect 2670 -2850 2740 -2780
rect 2780 -2850 2850 -2780
rect 2890 -2850 2960 -2780
rect 3000 -2850 3070 -2780
rect 1570 -2960 1640 -2890
rect 1680 -2960 1750 -2890
rect 1790 -2960 1860 -2890
rect 1900 -2960 1970 -2890
rect 2010 -2960 2080 -2890
rect 2120 -2960 2190 -2890
rect 2230 -2960 2300 -2890
rect 2340 -2960 2410 -2890
rect 2450 -2960 2520 -2890
rect 2560 -2960 2630 -2890
rect 2670 -2960 2740 -2890
rect 2780 -2960 2850 -2890
rect 2890 -2960 2960 -2890
rect 3000 -2960 3070 -2890
rect 11790 -2850 11860 -2780
rect 11900 -2850 11970 -2780
rect 12010 -2850 12080 -2780
rect 12120 -2850 12190 -2780
rect 12230 -2850 12300 -2780
rect 12340 -2850 12410 -2780
rect 12450 -2850 12520 -2780
rect 12560 -2850 12630 -2780
rect 12670 -2850 12740 -2780
rect 12780 -2850 12850 -2780
rect 12890 -2850 12960 -2780
rect 13000 -2850 13070 -2780
rect 13110 -2850 13180 -2780
rect 13220 -2850 13290 -2780
rect 11790 -2960 11860 -2890
rect 11900 -2960 11970 -2890
rect 12010 -2960 12080 -2890
rect 12120 -2960 12190 -2890
rect 12230 -2960 12300 -2890
rect 12340 -2960 12410 -2890
rect 12450 -2960 12520 -2890
rect 12560 -2960 12630 -2890
rect 12670 -2960 12740 -2890
rect 12780 -2960 12850 -2890
rect 12890 -2960 12960 -2890
rect 13000 -2960 13070 -2890
rect 13110 -2960 13180 -2890
rect 13220 -2960 13290 -2890
rect 22340 -3120 22410 -3050
rect 22450 -3120 22520 -3050
rect 22560 -3120 22630 -3050
rect 22340 -3230 22410 -3160
rect 22450 -3230 22520 -3160
rect 22560 -3230 22630 -3160
rect 22340 -3340 22410 -3270
rect 22450 -3340 22520 -3270
rect 22560 -3340 22630 -3270
rect 20070 -3760 20140 -3690
rect 20180 -3760 20250 -3690
rect 20290 -3760 20360 -3690
rect 20400 -3760 20470 -3690
rect 20070 -3870 20140 -3800
rect 20180 -3870 20250 -3800
rect 20290 -3870 20360 -3800
rect 20400 -3870 20470 -3800
rect 24550 -3760 24620 -3690
rect 24660 -3760 24730 -3690
rect 24770 -3760 24840 -3690
rect 24880 -3760 24950 -3690
rect 24550 -3870 24620 -3800
rect 24660 -3870 24730 -3800
rect 24770 -3870 24840 -3800
rect 24880 -3870 24950 -3800
rect -2200 -4540 -2130 -4470
rect -2090 -4540 -2020 -4470
rect -2200 -4650 -2130 -4580
rect -2090 -4650 -2020 -4580
rect -2200 -4760 -2130 -4690
rect -2090 -4760 -2020 -4690
rect -2200 -4870 -2130 -4800
rect -2090 -4870 -2020 -4800
rect 7310 -4630 7380 -4560
rect 7420 -4630 7490 -4560
rect 7530 -4630 7600 -4560
rect 7310 -4740 7380 -4670
rect 7420 -4740 7490 -4670
rect 7530 -4740 7600 -4670
rect 7310 -4850 7380 -4780
rect 7420 -4850 7490 -4780
rect 7530 -4850 7600 -4780
rect -2140 -5310 -2070 -5240
rect -2030 -5310 -1960 -5240
rect -2140 -5420 -2070 -5350
rect -2030 -5420 -1960 -5350
rect -2140 -5530 -2070 -5460
rect -2030 -5530 -1960 -5460
rect -2140 -5640 -2070 -5570
rect -2030 -5640 -1960 -5570
rect -840 -6570 -770 -6500
rect -710 -6570 -640 -6500
rect -840 -6680 -770 -6610
rect -710 -6680 -640 -6610
rect 7050 -6520 7110 -6460
rect 7150 -6520 7210 -6460
rect 7250 -6520 7310 -6460
rect 7050 -6620 7110 -6560
rect 7150 -6620 7210 -6560
rect 7250 -6620 7310 -6560
rect -840 -6790 -770 -6720
rect -710 -6790 -640 -6720
rect -840 -6900 -770 -6830
rect -710 -6900 -640 -6830
rect 4770 -6730 4830 -6670
rect 4870 -6730 4930 -6670
rect 4970 -6730 5030 -6670
rect 4770 -6830 4830 -6770
rect 4870 -6830 4930 -6770
rect 4970 -6830 5030 -6770
rect 7050 -6720 7110 -6660
rect 7150 -6720 7210 -6660
rect 7250 -6720 7310 -6660
rect 7050 -6820 7110 -6760
rect 7150 -6820 7210 -6760
rect 7250 -6820 7310 -6760
rect 7590 -6520 7650 -6460
rect 7690 -6520 7750 -6460
rect 7790 -6520 7850 -6460
rect 7590 -6620 7650 -6560
rect 7690 -6620 7750 -6560
rect 7790 -6620 7850 -6560
rect 15420 -6570 15490 -6500
rect 15550 -6570 15620 -6500
rect 7590 -6720 7650 -6660
rect 7690 -6720 7750 -6660
rect 7790 -6720 7850 -6660
rect 7590 -6820 7650 -6760
rect 7690 -6820 7750 -6760
rect 7790 -6820 7850 -6760
rect 9870 -6730 9930 -6670
rect 9970 -6730 10030 -6670
rect 10070 -6730 10130 -6670
rect 9870 -6830 9930 -6770
rect 9970 -6830 10030 -6770
rect 10070 -6830 10130 -6770
rect 4770 -6930 4830 -6870
rect 4870 -6930 4930 -6870
rect 4970 -6930 5030 -6870
rect 9870 -6930 9930 -6870
rect 9970 -6930 10030 -6870
rect 10070 -6930 10130 -6870
rect 15420 -6680 15490 -6610
rect 15550 -6680 15620 -6610
rect 15420 -6790 15490 -6720
rect 15550 -6790 15620 -6720
rect 15420 -6900 15490 -6830
rect 15550 -6900 15620 -6830
rect -2200 -7940 -2130 -7870
rect -2090 -7940 -2020 -7870
rect -2200 -8050 -2130 -7980
rect -2090 -8050 -2020 -7980
rect -2200 -8160 -2130 -8090
rect -2090 -8160 -2020 -8090
rect -2200 -8270 -2130 -8200
rect -2090 -8270 -2020 -8200
rect 14600 -8300 14670 -8230
rect 14700 -8300 14770 -8230
rect 14810 -8300 14880 -8230
rect 14600 -8410 14670 -8340
rect 14700 -8410 14770 -8340
rect 14810 -8410 14880 -8340
rect 14600 -8520 14670 -8450
rect 14700 -8520 14770 -8450
rect 14810 -8520 14880 -8450
rect -2140 -8710 -2070 -8640
rect -2030 -8710 -1960 -8640
rect -2140 -8820 -2070 -8750
rect -2030 -8820 -1960 -8750
rect -2140 -8930 -2070 -8860
rect -2030 -8930 -1960 -8860
rect -2140 -9040 -2070 -8970
rect -2030 -9040 -1960 -8970
rect 19230 -8630 19300 -8560
rect 19330 -8630 19400 -8560
rect 19430 -8630 19500 -8560
rect 19230 -8730 19300 -8660
rect 19330 -8730 19400 -8660
rect 19430 -8730 19500 -8660
rect 19230 -8830 19300 -8760
rect 19330 -8830 19400 -8760
rect 19430 -8830 19500 -8760
rect 19960 -9070 20030 -9000
rect 20060 -9070 20130 -9000
rect 20160 -9070 20230 -9000
rect 19960 -9170 20030 -9100
rect 20060 -9170 20130 -9100
rect 20160 -9170 20230 -9100
rect 19960 -9270 20030 -9200
rect 20060 -9270 20130 -9200
rect 20160 -9270 20230 -9200
rect -240 -9730 -170 -9660
rect -130 -9730 -60 -9660
rect -20 -9730 50 -9660
rect 90 -9730 160 -9660
rect -240 -9860 -170 -9790
rect -130 -9860 -60 -9790
rect -20 -9860 50 -9790
rect 90 -9860 160 -9790
rect 14720 -9730 14790 -9660
rect 14830 -9730 14900 -9660
rect 14940 -9730 15010 -9660
rect 15050 -9730 15120 -9660
rect 14720 -9860 14790 -9790
rect 14830 -9860 14900 -9790
rect 14940 -9860 15010 -9790
rect 15050 -9860 15120 -9790
rect 1150 -10410 1220 -10340
rect 1260 -10410 1330 -10340
rect 1370 -10410 1440 -10340
rect 1480 -10410 1550 -10340
rect 1590 -10410 1660 -10340
rect 1700 -10410 1770 -10340
rect 1810 -10410 1880 -10340
rect 1920 -10410 1990 -10340
rect 2030 -10410 2100 -10340
rect 2140 -10410 2210 -10340
rect 2250 -10410 2320 -10340
rect 2360 -10410 2430 -10340
rect 2470 -10410 2540 -10340
rect 2580 -10410 2650 -10340
rect 1150 -10520 1220 -10450
rect 1260 -10520 1330 -10450
rect 1370 -10520 1440 -10450
rect 1480 -10520 1550 -10450
rect 1590 -10520 1660 -10450
rect 1700 -10520 1770 -10450
rect 1810 -10520 1880 -10450
rect 1920 -10520 1990 -10450
rect 2030 -10520 2100 -10450
rect 2140 -10520 2210 -10450
rect 2250 -10520 2320 -10450
rect 2360 -10520 2430 -10450
rect 2470 -10520 2540 -10450
rect 2580 -10520 2650 -10450
rect 12290 -10440 12360 -10370
rect 12400 -10440 12470 -10370
rect 12510 -10440 12580 -10370
rect 12620 -10440 12690 -10370
rect 12730 -10440 12800 -10370
rect 12840 -10440 12910 -10370
rect 12950 -10440 13020 -10370
rect 13060 -10440 13130 -10370
rect 13170 -10440 13240 -10370
rect 13280 -10440 13350 -10370
rect 13390 -10440 13460 -10370
rect 13500 -10440 13570 -10370
rect 13610 -10440 13680 -10370
rect 13720 -10440 13790 -10370
rect 12290 -10550 12360 -10480
rect 12400 -10550 12470 -10480
rect 12510 -10550 12580 -10480
rect 12620 -10550 12690 -10480
rect 12730 -10550 12800 -10480
rect 12840 -10550 12910 -10480
rect 12950 -10550 13020 -10480
rect 13060 -10550 13130 -10480
rect 13170 -10550 13240 -10480
rect 13280 -10550 13350 -10480
rect 13390 -10550 13460 -10480
rect 13500 -10550 13570 -10480
rect 13610 -10550 13680 -10480
rect 13720 -10550 13790 -10480
rect 2240 -12370 2310 -12300
rect 2350 -12370 2420 -12300
rect 2460 -12370 2530 -12300
rect 2570 -12370 2640 -12300
rect 2680 -12370 2750 -12300
rect 2790 -12370 2860 -12300
rect 2900 -12370 2970 -12300
rect 3010 -12370 3080 -12300
rect 3120 -12370 3190 -12300
rect 3230 -12370 3300 -12300
rect 3340 -12370 3410 -12300
rect 3450 -12370 3520 -12300
rect 3560 -12370 3630 -12300
rect 3670 -12370 3740 -12300
rect 2240 -12480 2310 -12410
rect 2350 -12480 2420 -12410
rect 2460 -12480 2530 -12410
rect 2570 -12480 2640 -12410
rect 2680 -12480 2750 -12410
rect 2790 -12480 2860 -12410
rect 2900 -12480 2970 -12410
rect 3010 -12480 3080 -12410
rect 3120 -12480 3190 -12410
rect 3230 -12480 3300 -12410
rect 3340 -12480 3410 -12410
rect 3450 -12480 3520 -12410
rect 3560 -12480 3630 -12410
rect 3670 -12480 3740 -12410
rect 11120 -12370 11190 -12300
rect 11230 -12370 11300 -12300
rect 11340 -12370 11410 -12300
rect 11450 -12370 11520 -12300
rect 11560 -12370 11630 -12300
rect 11670 -12370 11740 -12300
rect 11780 -12370 11850 -12300
rect 11890 -12370 11960 -12300
rect 12000 -12370 12070 -12300
rect 12110 -12370 12180 -12300
rect 12220 -12370 12290 -12300
rect 12330 -12370 12400 -12300
rect 12440 -12370 12510 -12300
rect 12550 -12370 12620 -12300
rect 11120 -12480 11190 -12410
rect 11230 -12480 11300 -12410
rect 11340 -12480 11410 -12410
rect 11450 -12480 11520 -12410
rect 11560 -12480 11630 -12410
rect 11670 -12480 11740 -12410
rect 11780 -12480 11850 -12410
rect 11890 -12480 11960 -12410
rect 12000 -12480 12070 -12410
rect 12110 -12480 12180 -12410
rect 12220 -12480 12290 -12410
rect 12330 -12480 12400 -12410
rect 12440 -12480 12510 -12410
rect 12550 -12480 12620 -12410
rect 7010 -13310 7070 -13250
rect 7110 -13310 7170 -13250
rect 7210 -13310 7270 -13250
rect 7010 -13400 7070 -13340
rect 7110 -13400 7170 -13340
rect 7210 -13400 7270 -13340
rect 7010 -13490 7070 -13430
rect 7110 -13490 7170 -13430
rect 7210 -13490 7270 -13430
rect 7010 -13590 7070 -13530
rect 7110 -13590 7170 -13530
rect 7210 -13590 7270 -13530
rect 7010 -13680 7070 -13620
rect 7110 -13680 7170 -13620
rect 7210 -13680 7270 -13620
rect 7010 -13770 7070 -13710
rect 7110 -13770 7170 -13710
rect 7210 -13770 7270 -13710
rect 7630 -13310 7690 -13250
rect 7730 -13310 7790 -13250
rect 7830 -13310 7890 -13250
rect 7630 -13400 7690 -13340
rect 7730 -13400 7790 -13340
rect 7830 -13400 7890 -13340
rect 7630 -13490 7690 -13430
rect 7730 -13490 7790 -13430
rect 7830 -13490 7890 -13430
rect 7630 -13590 7690 -13530
rect 7730 -13590 7790 -13530
rect 7830 -13590 7890 -13530
rect 7630 -13680 7690 -13620
rect 7730 -13680 7790 -13620
rect 7830 -13680 7890 -13620
rect 7630 -13770 7690 -13710
rect 7730 -13770 7790 -13710
rect 7830 -13770 7890 -13710
rect 19230 -14290 19300 -14220
rect 19330 -14290 19400 -14220
rect 19430 -14290 19500 -14220
rect 19230 -14390 19300 -14320
rect 19330 -14390 19400 -14320
rect 19430 -14390 19500 -14320
rect 19230 -14490 19300 -14420
rect 19330 -14490 19400 -14420
rect 19430 -14490 19500 -14420
rect 20480 -14940 20550 -14870
rect 20580 -14940 20650 -14870
rect 20680 -14940 20750 -14870
rect 20480 -15040 20550 -14970
rect 20580 -15040 20650 -14970
rect 20680 -15040 20750 -14970
rect 20480 -15140 20550 -15070
rect 20580 -15140 20650 -15070
rect 20680 -15140 20750 -15070
rect 5040 -17160 5100 -17100
rect 5140 -17160 5200 -17100
rect 5240 -17160 5300 -17100
rect 5040 -17260 5100 -17200
rect 5140 -17260 5200 -17200
rect 5240 -17260 5300 -17200
rect 5040 -17360 5100 -17300
rect 5140 -17360 5200 -17300
rect 5240 -17360 5300 -17300
rect 9600 -17160 9660 -17100
rect 9700 -17160 9760 -17100
rect 9800 -17160 9860 -17100
rect 9600 -17260 9660 -17200
rect 9700 -17260 9760 -17200
rect 9800 -17260 9860 -17200
rect 9600 -17360 9660 -17300
rect 9700 -17360 9760 -17300
rect 9800 -17360 9860 -17300
rect 7230 -17670 7300 -17600
rect 7340 -17670 7410 -17600
rect 7450 -17670 7520 -17600
rect 7560 -17670 7630 -17600
rect 7230 -17780 7300 -17710
rect 7340 -17780 7410 -17710
rect 7450 -17780 7520 -17710
rect 7560 -17780 7630 -17710
rect 7230 -17890 7300 -17820
rect 7340 -17890 7410 -17820
rect 7450 -17890 7520 -17820
rect 7560 -17890 7630 -17820
rect 7230 -18000 7300 -17930
rect 7340 -18000 7410 -17930
rect 7450 -18000 7520 -17930
rect 7560 -18000 7630 -17930
rect 19230 -20360 19300 -20290
rect 19330 -20360 19400 -20290
rect 19430 -20360 19500 -20290
rect 19230 -20460 19300 -20390
rect 19330 -20460 19400 -20390
rect 19430 -20460 19500 -20390
rect 19230 -20560 19300 -20490
rect 19330 -20560 19400 -20490
rect 19430 -20560 19500 -20490
rect 20040 -20790 20110 -20720
rect 20140 -20790 20210 -20720
rect 20240 -20790 20310 -20720
rect 20040 -20890 20110 -20820
rect 20140 -20890 20210 -20820
rect 20240 -20890 20310 -20820
rect 20040 -20990 20110 -20920
rect 20140 -20990 20210 -20920
rect 20240 -20990 20310 -20920
rect 2280 -22730 2350 -22660
rect 2390 -22730 2460 -22660
rect 2500 -22730 2570 -22660
rect 2610 -22730 2680 -22660
rect 2720 -22730 2790 -22660
rect 2830 -22730 2900 -22660
rect 2940 -22730 3010 -22660
rect 3050 -22730 3120 -22660
rect 3160 -22730 3230 -22660
rect 3270 -22730 3340 -22660
rect 3380 -22730 3450 -22660
rect 3490 -22730 3560 -22660
rect 3600 -22730 3670 -22660
rect 3710 -22730 3780 -22660
rect 2280 -22840 2350 -22770
rect 2390 -22840 2460 -22770
rect 2500 -22840 2570 -22770
rect 2610 -22840 2680 -22770
rect 2720 -22840 2790 -22770
rect 2830 -22840 2900 -22770
rect 2940 -22840 3010 -22770
rect 3050 -22840 3120 -22770
rect 3160 -22840 3230 -22770
rect 3270 -22840 3340 -22770
rect 3380 -22840 3450 -22770
rect 3490 -22840 3560 -22770
rect 3600 -22840 3670 -22770
rect 3710 -22840 3780 -22770
rect 11160 -22730 11230 -22660
rect 11270 -22730 11340 -22660
rect 11380 -22730 11450 -22660
rect 11490 -22730 11560 -22660
rect 11600 -22730 11670 -22660
rect 11710 -22730 11780 -22660
rect 11820 -22730 11890 -22660
rect 11930 -22730 12000 -22660
rect 12040 -22730 12110 -22660
rect 12150 -22730 12220 -22660
rect 12260 -22730 12330 -22660
rect 12370 -22730 12440 -22660
rect 12480 -22730 12550 -22660
rect 12590 -22730 12660 -22660
rect 11160 -22840 11230 -22770
rect 11270 -22840 11340 -22770
rect 11380 -22840 11450 -22770
rect 11490 -22840 11560 -22770
rect 11600 -22840 11670 -22770
rect 11710 -22840 11780 -22770
rect 11820 -22840 11890 -22770
rect 11930 -22840 12000 -22770
rect 12040 -22840 12110 -22770
rect 12150 -22840 12220 -22770
rect 12260 -22840 12330 -22770
rect 12370 -22840 12440 -22770
rect 12480 -22840 12550 -22770
rect 12590 -22840 12660 -22770
<< metal3 >>
rect -5020 8500 7290 21140
rect -5020 8430 -4730 8500
rect -4660 8430 -4640 8500
rect -4570 8430 -4550 8500
rect -4480 8430 -4460 8500
rect -4390 8430 -4370 8500
rect -4300 8430 -4280 8500
rect -4210 8430 -4190 8500
rect -4120 8430 -4100 8500
rect -4030 8430 -4010 8500
rect -3940 8430 -3920 8500
rect -3850 8430 -3830 8500
rect -3760 8430 -3740 8500
rect -3670 8430 -3650 8500
rect -3580 8430 -3560 8500
rect -3490 8430 -3470 8500
rect -3400 8430 -3380 8500
rect -3310 8430 -3290 8500
rect -3220 8430 -3200 8500
rect -3130 8430 -3110 8500
rect -3040 8430 -3020 8500
rect -2950 8430 -2930 8500
rect -2860 8430 -2840 8500
rect -2770 8430 -2750 8500
rect -2680 8430 -2660 8500
rect -2590 8430 -2570 8500
rect -2500 8430 -2480 8500
rect -2410 8430 -2390 8500
rect -2320 8430 -2300 8500
rect -2230 8430 -2210 8500
rect -2140 8430 -2120 8500
rect -2050 8430 -2030 8500
rect -1960 8430 -1940 8500
rect -1870 8430 -1850 8500
rect -1780 8430 -1720 8500
rect -1650 8430 -1630 8500
rect -1560 8430 -1540 8500
rect -1470 8430 -1450 8500
rect -1380 8430 -1360 8500
rect -1290 8430 -1270 8500
rect -1200 8430 -1180 8500
rect -1110 8430 -1090 8500
rect -1020 8430 -1000 8500
rect -930 8430 -910 8500
rect -840 8430 -820 8500
rect -750 8430 -730 8500
rect -660 8430 -640 8500
rect -570 8430 -550 8500
rect -480 8430 -460 8500
rect -390 8430 -370 8500
rect -300 8430 -280 8500
rect -210 8430 -190 8500
rect -120 8430 -100 8500
rect -30 8430 -10 8500
rect 60 8430 80 8500
rect 150 8430 170 8500
rect 240 8430 260 8500
rect 330 8430 350 8500
rect 420 8430 440 8500
rect 510 8430 530 8500
rect 600 8430 620 8500
rect 690 8430 710 8500
rect 780 8430 800 8500
rect 870 8430 890 8500
rect 960 8430 980 8500
rect 1050 8430 1070 8500
rect 1140 8430 1160 8500
rect 1230 8430 1290 8500
rect 1360 8430 1380 8500
rect 1450 8430 1470 8500
rect 1540 8430 1560 8500
rect 1630 8430 1650 8500
rect 1720 8430 1740 8500
rect 1810 8430 1830 8500
rect 1900 8430 1920 8500
rect 1990 8430 2010 8500
rect 2080 8430 2100 8500
rect 2170 8430 2190 8500
rect 2260 8430 2280 8500
rect 2350 8430 2370 8500
rect 2440 8430 2460 8500
rect 2530 8430 2550 8500
rect 2620 8430 2640 8500
rect 2710 8430 2730 8500
rect 2800 8430 2820 8500
rect 2890 8430 2910 8500
rect 2980 8430 3000 8500
rect 3070 8430 3090 8500
rect 3160 8430 3180 8500
rect 3250 8430 3270 8500
rect 3340 8430 3360 8500
rect 3430 8430 3450 8500
rect 3520 8430 3540 8500
rect 3610 8430 3630 8500
rect 3700 8430 3720 8500
rect 3790 8430 3810 8500
rect 3880 8430 3900 8500
rect 3970 8430 3990 8500
rect 4060 8430 4080 8500
rect 4150 8430 4170 8500
rect 4240 8430 4300 8500
rect 4370 8430 4390 8500
rect 4460 8430 4480 8500
rect 4550 8430 4570 8500
rect 4640 8430 4660 8500
rect 4730 8430 4750 8500
rect 4820 8430 4840 8500
rect 4910 8430 4930 8500
rect 5000 8430 5020 8500
rect 5090 8430 5110 8500
rect 5180 8430 5200 8500
rect 5270 8430 5290 8500
rect 5360 8430 5380 8500
rect 5450 8430 5470 8500
rect 5540 8430 5560 8500
rect 5630 8430 5650 8500
rect 5720 8430 5740 8500
rect 5810 8430 5830 8500
rect 5900 8430 5920 8500
rect 5990 8430 6010 8500
rect 6080 8430 6100 8500
rect 6170 8430 6190 8500
rect 6260 8430 6280 8500
rect 6350 8430 6370 8500
rect 6440 8430 6460 8500
rect 6530 8430 6550 8500
rect 6620 8430 6640 8500
rect 6710 8430 6730 8500
rect 6800 8430 6820 8500
rect 6890 8430 6910 8500
rect 6980 8430 7000 8500
rect 7070 8430 7090 8500
rect 7160 8430 7180 8500
rect 7250 8430 7290 8500
rect -5020 8410 7290 8430
rect -5020 8340 -4730 8410
rect -4660 8340 -4640 8410
rect -4570 8340 -4550 8410
rect -4480 8340 -4460 8410
rect -4390 8340 -4370 8410
rect -4300 8340 -4280 8410
rect -4210 8340 -4190 8410
rect -4120 8340 -4100 8410
rect -4030 8340 -4010 8410
rect -3940 8340 -3920 8410
rect -3850 8340 -3830 8410
rect -3760 8340 -3740 8410
rect -3670 8340 -3650 8410
rect -3580 8340 -3560 8410
rect -3490 8340 -3470 8410
rect -3400 8340 -3380 8410
rect -3310 8340 -3290 8410
rect -3220 8340 -3200 8410
rect -3130 8340 -3110 8410
rect -3040 8340 -3020 8410
rect -2950 8340 -2930 8410
rect -2860 8340 -2840 8410
rect -2770 8340 -2750 8410
rect -2680 8340 -2660 8410
rect -2590 8340 -2570 8410
rect -2500 8340 -2480 8410
rect -2410 8340 -2390 8410
rect -2320 8340 -2300 8410
rect -2230 8340 -2210 8410
rect -2140 8340 -2120 8410
rect -2050 8340 -2030 8410
rect -1960 8340 -1940 8410
rect -1870 8340 -1850 8410
rect -1780 8340 -1720 8410
rect -1650 8340 -1630 8410
rect -1560 8340 -1540 8410
rect -1470 8340 -1450 8410
rect -1380 8340 -1360 8410
rect -1290 8340 -1270 8410
rect -1200 8340 -1180 8410
rect -1110 8340 -1090 8410
rect -1020 8340 -1000 8410
rect -930 8340 -910 8410
rect -840 8340 -820 8410
rect -750 8340 -730 8410
rect -660 8340 -640 8410
rect -570 8340 -550 8410
rect -480 8340 -460 8410
rect -390 8340 -370 8410
rect -300 8340 -280 8410
rect -210 8340 -190 8410
rect -120 8340 -100 8410
rect -30 8340 -10 8410
rect 60 8340 80 8410
rect 150 8340 170 8410
rect 240 8340 260 8410
rect 330 8340 350 8410
rect 420 8340 440 8410
rect 510 8340 530 8410
rect 600 8340 620 8410
rect 690 8340 710 8410
rect 780 8340 800 8410
rect 870 8340 890 8410
rect 960 8340 980 8410
rect 1050 8340 1070 8410
rect 1140 8340 1160 8410
rect 1230 8340 1290 8410
rect 1360 8340 1380 8410
rect 1450 8340 1470 8410
rect 1540 8340 1560 8410
rect 1630 8340 1650 8410
rect 1720 8340 1740 8410
rect 1810 8340 1830 8410
rect 1900 8340 1920 8410
rect 1990 8340 2010 8410
rect 2080 8340 2100 8410
rect 2170 8340 2190 8410
rect 2260 8340 2280 8410
rect 2350 8340 2370 8410
rect 2440 8340 2460 8410
rect 2530 8340 2550 8410
rect 2620 8340 2640 8410
rect 2710 8340 2730 8410
rect 2800 8340 2820 8410
rect 2890 8340 2910 8410
rect 2980 8340 3000 8410
rect 3070 8340 3090 8410
rect 3160 8340 3180 8410
rect 3250 8340 3270 8410
rect 3340 8340 3360 8410
rect 3430 8340 3450 8410
rect 3520 8340 3540 8410
rect 3610 8340 3630 8410
rect 3700 8340 3720 8410
rect 3790 8340 3810 8410
rect 3880 8340 3900 8410
rect 3970 8340 3990 8410
rect 4060 8340 4080 8410
rect 4150 8340 4170 8410
rect 4240 8340 4300 8410
rect 4370 8340 4390 8410
rect 4460 8340 4480 8410
rect 4550 8340 4570 8410
rect 4640 8340 4660 8410
rect 4730 8340 4750 8410
rect 4820 8340 4840 8410
rect 4910 8340 4930 8410
rect 5000 8340 5020 8410
rect 5090 8340 5110 8410
rect 5180 8340 5200 8410
rect 5270 8340 5290 8410
rect 5360 8340 5380 8410
rect 5450 8340 5470 8410
rect 5540 8340 5560 8410
rect 5630 8340 5650 8410
rect 5720 8340 5740 8410
rect 5810 8340 5830 8410
rect 5900 8340 5920 8410
rect 5990 8340 6010 8410
rect 6080 8340 6100 8410
rect 6170 8340 6190 8410
rect 6260 8340 6280 8410
rect 6350 8340 6370 8410
rect 6440 8340 6460 8410
rect 6530 8340 6550 8410
rect 6620 8340 6640 8410
rect 6710 8340 6730 8410
rect 6800 8340 6820 8410
rect 6890 8340 6910 8410
rect 6980 8340 7000 8410
rect 7070 8340 7090 8410
rect 7160 8340 7180 8410
rect 7250 8340 7290 8410
rect -5020 8320 7290 8340
rect -5020 8250 -4730 8320
rect -4660 8250 -4640 8320
rect -4570 8250 -4550 8320
rect -4480 8250 -4460 8320
rect -4390 8250 -4370 8320
rect -4300 8250 -4280 8320
rect -4210 8250 -4190 8320
rect -4120 8250 -4100 8320
rect -4030 8250 -4010 8320
rect -3940 8250 -3920 8320
rect -3850 8250 -3830 8320
rect -3760 8250 -3740 8320
rect -3670 8250 -3650 8320
rect -3580 8250 -3560 8320
rect -3490 8250 -3470 8320
rect -3400 8250 -3380 8320
rect -3310 8250 -3290 8320
rect -3220 8250 -3200 8320
rect -3130 8250 -3110 8320
rect -3040 8250 -3020 8320
rect -2950 8250 -2930 8320
rect -2860 8250 -2840 8320
rect -2770 8250 -2750 8320
rect -2680 8250 -2660 8320
rect -2590 8250 -2570 8320
rect -2500 8250 -2480 8320
rect -2410 8250 -2390 8320
rect -2320 8250 -2300 8320
rect -2230 8250 -2210 8320
rect -2140 8250 -2120 8320
rect -2050 8250 -2030 8320
rect -1960 8250 -1940 8320
rect -1870 8250 -1850 8320
rect -1780 8250 -1720 8320
rect -1650 8250 -1630 8320
rect -1560 8250 -1540 8320
rect -1470 8250 -1450 8320
rect -1380 8250 -1360 8320
rect -1290 8250 -1270 8320
rect -1200 8250 -1180 8320
rect -1110 8250 -1090 8320
rect -1020 8250 -1000 8320
rect -930 8250 -910 8320
rect -840 8250 -820 8320
rect -750 8250 -730 8320
rect -660 8250 -640 8320
rect -570 8250 -550 8320
rect -480 8250 -460 8320
rect -390 8250 -370 8320
rect -300 8250 -280 8320
rect -210 8250 -190 8320
rect -120 8250 -100 8320
rect -30 8250 -10 8320
rect 60 8250 80 8320
rect 150 8250 170 8320
rect 240 8250 260 8320
rect 330 8250 350 8320
rect 420 8250 440 8320
rect 510 8250 530 8320
rect 600 8250 620 8320
rect 690 8250 710 8320
rect 780 8250 800 8320
rect 870 8250 890 8320
rect 960 8250 980 8320
rect 1050 8250 1070 8320
rect 1140 8250 1160 8320
rect 1230 8250 1290 8320
rect 1360 8250 1380 8320
rect 1450 8250 1470 8320
rect 1540 8250 1560 8320
rect 1630 8250 1650 8320
rect 1720 8250 1740 8320
rect 1810 8250 1830 8320
rect 1900 8250 1920 8320
rect 1990 8250 2010 8320
rect 2080 8250 2100 8320
rect 2170 8250 2190 8320
rect 2260 8250 2280 8320
rect 2350 8250 2370 8320
rect 2440 8250 2460 8320
rect 2530 8250 2550 8320
rect 2620 8250 2640 8320
rect 2710 8250 2730 8320
rect 2800 8250 2820 8320
rect 2890 8250 2910 8320
rect 2980 8250 3000 8320
rect 3070 8250 3090 8320
rect 3160 8250 3180 8320
rect 3250 8250 3270 8320
rect 3340 8250 3360 8320
rect 3430 8250 3450 8320
rect 3520 8250 3540 8320
rect 3610 8250 3630 8320
rect 3700 8250 3720 8320
rect 3790 8250 3810 8320
rect 3880 8250 3900 8320
rect 3970 8250 3990 8320
rect 4060 8250 4080 8320
rect 4150 8250 4170 8320
rect 4240 8250 4300 8320
rect 4370 8250 4390 8320
rect 4460 8250 4480 8320
rect 4550 8250 4570 8320
rect 4640 8250 4660 8320
rect 4730 8250 4750 8320
rect 4820 8250 4840 8320
rect 4910 8250 4930 8320
rect 5000 8250 5020 8320
rect 5090 8250 5110 8320
rect 5180 8250 5200 8320
rect 5270 8250 5290 8320
rect 5360 8250 5380 8320
rect 5450 8250 5470 8320
rect 5540 8250 5560 8320
rect 5630 8250 5650 8320
rect 5720 8250 5740 8320
rect 5810 8250 5830 8320
rect 5900 8250 5920 8320
rect 5990 8250 6010 8320
rect 6080 8250 6100 8320
rect 6170 8250 6190 8320
rect 6260 8250 6280 8320
rect 6350 8250 6370 8320
rect 6440 8250 6460 8320
rect 6530 8250 6550 8320
rect 6620 8250 6640 8320
rect 6710 8250 6730 8320
rect 6800 8250 6820 8320
rect 6890 8250 6910 8320
rect 6980 8250 7000 8320
rect 7070 8250 7090 8320
rect 7160 8250 7180 8320
rect 7250 8250 7290 8320
rect -5020 8190 7290 8250
rect 7610 8500 19920 21140
rect 7610 8430 7650 8500
rect 7720 8430 7740 8500
rect 7810 8430 7830 8500
rect 7900 8430 7920 8500
rect 7990 8430 8010 8500
rect 8080 8430 8100 8500
rect 8170 8430 8190 8500
rect 8260 8430 8280 8500
rect 8350 8430 8370 8500
rect 8440 8430 8460 8500
rect 8530 8430 8550 8500
rect 8620 8430 8640 8500
rect 8710 8430 8730 8500
rect 8800 8430 8820 8500
rect 8890 8430 8910 8500
rect 8980 8430 9000 8500
rect 9070 8430 9090 8500
rect 9160 8430 9180 8500
rect 9250 8430 9270 8500
rect 9340 8430 9360 8500
rect 9430 8430 9450 8500
rect 9520 8430 9540 8500
rect 9610 8430 9630 8500
rect 9700 8430 9720 8500
rect 9790 8430 9810 8500
rect 9880 8430 9900 8500
rect 9970 8430 9990 8500
rect 10060 8430 10080 8500
rect 10150 8430 10170 8500
rect 10240 8430 10260 8500
rect 10330 8430 10350 8500
rect 10420 8430 10440 8500
rect 10510 8430 10530 8500
rect 10600 8430 10660 8500
rect 10730 8430 10750 8500
rect 10820 8430 10840 8500
rect 10910 8430 10930 8500
rect 11000 8430 11020 8500
rect 11090 8430 11110 8500
rect 11180 8430 11200 8500
rect 11270 8430 11290 8500
rect 11360 8430 11380 8500
rect 11450 8430 11470 8500
rect 11540 8430 11560 8500
rect 11630 8430 11650 8500
rect 11720 8430 11740 8500
rect 11810 8430 11830 8500
rect 11900 8430 11920 8500
rect 11990 8430 12010 8500
rect 12080 8430 12100 8500
rect 12170 8430 12190 8500
rect 12260 8430 12280 8500
rect 12350 8430 12370 8500
rect 12440 8430 12460 8500
rect 12530 8430 12550 8500
rect 12620 8430 12640 8500
rect 12710 8430 12730 8500
rect 12800 8430 12820 8500
rect 12890 8430 12910 8500
rect 12980 8430 13000 8500
rect 13070 8430 13090 8500
rect 13160 8430 13180 8500
rect 13250 8430 13270 8500
rect 13340 8430 13360 8500
rect 13430 8430 13450 8500
rect 13520 8430 13540 8500
rect 13610 8430 13670 8500
rect 13740 8430 13760 8500
rect 13830 8430 13850 8500
rect 13920 8430 13940 8500
rect 14010 8430 14030 8500
rect 14100 8430 14120 8500
rect 14190 8430 14210 8500
rect 14280 8430 14300 8500
rect 14370 8430 14390 8500
rect 14460 8430 14480 8500
rect 14550 8430 14570 8500
rect 14640 8430 14660 8500
rect 14730 8430 14750 8500
rect 14820 8430 14840 8500
rect 14910 8430 14930 8500
rect 15000 8430 15020 8500
rect 15090 8430 15110 8500
rect 15180 8430 15200 8500
rect 15270 8430 15290 8500
rect 15360 8430 15380 8500
rect 15450 8430 15470 8500
rect 15540 8430 15560 8500
rect 15630 8430 15650 8500
rect 15720 8430 15740 8500
rect 15810 8430 15830 8500
rect 15900 8430 15920 8500
rect 15990 8430 16010 8500
rect 16080 8430 16100 8500
rect 16170 8430 16190 8500
rect 16260 8430 16280 8500
rect 16350 8430 16370 8500
rect 16440 8430 16460 8500
rect 16530 8430 16550 8500
rect 16620 8430 16680 8500
rect 16750 8430 16770 8500
rect 16840 8430 16860 8500
rect 16930 8430 16950 8500
rect 17020 8430 17040 8500
rect 17110 8430 17130 8500
rect 17200 8430 17220 8500
rect 17290 8430 17310 8500
rect 17380 8430 17400 8500
rect 17470 8430 17490 8500
rect 17560 8430 17580 8500
rect 17650 8430 17670 8500
rect 17740 8430 17760 8500
rect 17830 8430 17850 8500
rect 17920 8430 17940 8500
rect 18010 8430 18030 8500
rect 18100 8430 18120 8500
rect 18190 8430 18210 8500
rect 18280 8430 18300 8500
rect 18370 8430 18390 8500
rect 18460 8430 18480 8500
rect 18550 8430 18570 8500
rect 18640 8430 18660 8500
rect 18730 8430 18750 8500
rect 18820 8430 18840 8500
rect 18910 8430 18930 8500
rect 19000 8430 19020 8500
rect 19090 8430 19110 8500
rect 19180 8430 19200 8500
rect 19270 8430 19290 8500
rect 19360 8430 19380 8500
rect 19450 8430 19470 8500
rect 19540 8430 19560 8500
rect 19630 8430 19920 8500
rect 7610 8410 19920 8430
rect 7610 8340 7650 8410
rect 7720 8340 7740 8410
rect 7810 8340 7830 8410
rect 7900 8340 7920 8410
rect 7990 8340 8010 8410
rect 8080 8340 8100 8410
rect 8170 8340 8190 8410
rect 8260 8340 8280 8410
rect 8350 8340 8370 8410
rect 8440 8340 8460 8410
rect 8530 8340 8550 8410
rect 8620 8340 8640 8410
rect 8710 8340 8730 8410
rect 8800 8340 8820 8410
rect 8890 8340 8910 8410
rect 8980 8340 9000 8410
rect 9070 8340 9090 8410
rect 9160 8340 9180 8410
rect 9250 8340 9270 8410
rect 9340 8340 9360 8410
rect 9430 8340 9450 8410
rect 9520 8340 9540 8410
rect 9610 8340 9630 8410
rect 9700 8340 9720 8410
rect 9790 8340 9810 8410
rect 9880 8340 9900 8410
rect 9970 8340 9990 8410
rect 10060 8340 10080 8410
rect 10150 8340 10170 8410
rect 10240 8340 10260 8410
rect 10330 8340 10350 8410
rect 10420 8340 10440 8410
rect 10510 8340 10530 8410
rect 10600 8340 10660 8410
rect 10730 8340 10750 8410
rect 10820 8340 10840 8410
rect 10910 8340 10930 8410
rect 11000 8340 11020 8410
rect 11090 8340 11110 8410
rect 11180 8340 11200 8410
rect 11270 8340 11290 8410
rect 11360 8340 11380 8410
rect 11450 8340 11470 8410
rect 11540 8340 11560 8410
rect 11630 8340 11650 8410
rect 11720 8340 11740 8410
rect 11810 8340 11830 8410
rect 11900 8340 11920 8410
rect 11990 8340 12010 8410
rect 12080 8340 12100 8410
rect 12170 8340 12190 8410
rect 12260 8340 12280 8410
rect 12350 8340 12370 8410
rect 12440 8340 12460 8410
rect 12530 8340 12550 8410
rect 12620 8340 12640 8410
rect 12710 8340 12730 8410
rect 12800 8340 12820 8410
rect 12890 8340 12910 8410
rect 12980 8340 13000 8410
rect 13070 8340 13090 8410
rect 13160 8340 13180 8410
rect 13250 8340 13270 8410
rect 13340 8340 13360 8410
rect 13430 8340 13450 8410
rect 13520 8340 13540 8410
rect 13610 8340 13670 8410
rect 13740 8340 13760 8410
rect 13830 8340 13850 8410
rect 13920 8340 13940 8410
rect 14010 8340 14030 8410
rect 14100 8340 14120 8410
rect 14190 8340 14210 8410
rect 14280 8340 14300 8410
rect 14370 8340 14390 8410
rect 14460 8340 14480 8410
rect 14550 8340 14570 8410
rect 14640 8340 14660 8410
rect 14730 8340 14750 8410
rect 14820 8340 14840 8410
rect 14910 8340 14930 8410
rect 15000 8340 15020 8410
rect 15090 8340 15110 8410
rect 15180 8340 15200 8410
rect 15270 8340 15290 8410
rect 15360 8340 15380 8410
rect 15450 8340 15470 8410
rect 15540 8340 15560 8410
rect 15630 8340 15650 8410
rect 15720 8340 15740 8410
rect 15810 8340 15830 8410
rect 15900 8340 15920 8410
rect 15990 8340 16010 8410
rect 16080 8340 16100 8410
rect 16170 8340 16190 8410
rect 16260 8340 16280 8410
rect 16350 8340 16370 8410
rect 16440 8340 16460 8410
rect 16530 8340 16550 8410
rect 16620 8340 16680 8410
rect 16750 8340 16770 8410
rect 16840 8340 16860 8410
rect 16930 8340 16950 8410
rect 17020 8340 17040 8410
rect 17110 8340 17130 8410
rect 17200 8340 17220 8410
rect 17290 8340 17310 8410
rect 17380 8340 17400 8410
rect 17470 8340 17490 8410
rect 17560 8340 17580 8410
rect 17650 8340 17670 8410
rect 17740 8340 17760 8410
rect 17830 8340 17850 8410
rect 17920 8340 17940 8410
rect 18010 8340 18030 8410
rect 18100 8340 18120 8410
rect 18190 8340 18210 8410
rect 18280 8340 18300 8410
rect 18370 8340 18390 8410
rect 18460 8340 18480 8410
rect 18550 8340 18570 8410
rect 18640 8340 18660 8410
rect 18730 8340 18750 8410
rect 18820 8340 18840 8410
rect 18910 8340 18930 8410
rect 19000 8340 19020 8410
rect 19090 8340 19110 8410
rect 19180 8340 19200 8410
rect 19270 8340 19290 8410
rect 19360 8340 19380 8410
rect 19450 8340 19470 8410
rect 19540 8340 19560 8410
rect 19630 8340 19920 8410
rect 7610 8320 19920 8340
rect 7610 8250 7650 8320
rect 7720 8250 7740 8320
rect 7810 8250 7830 8320
rect 7900 8250 7920 8320
rect 7990 8250 8010 8320
rect 8080 8250 8100 8320
rect 8170 8250 8190 8320
rect 8260 8250 8280 8320
rect 8350 8250 8370 8320
rect 8440 8250 8460 8320
rect 8530 8250 8550 8320
rect 8620 8250 8640 8320
rect 8710 8250 8730 8320
rect 8800 8250 8820 8320
rect 8890 8250 8910 8320
rect 8980 8250 9000 8320
rect 9070 8250 9090 8320
rect 9160 8250 9180 8320
rect 9250 8250 9270 8320
rect 9340 8250 9360 8320
rect 9430 8250 9450 8320
rect 9520 8250 9540 8320
rect 9610 8250 9630 8320
rect 9700 8250 9720 8320
rect 9790 8250 9810 8320
rect 9880 8250 9900 8320
rect 9970 8250 9990 8320
rect 10060 8250 10080 8320
rect 10150 8250 10170 8320
rect 10240 8250 10260 8320
rect 10330 8250 10350 8320
rect 10420 8250 10440 8320
rect 10510 8250 10530 8320
rect 10600 8250 10660 8320
rect 10730 8250 10750 8320
rect 10820 8250 10840 8320
rect 10910 8250 10930 8320
rect 11000 8250 11020 8320
rect 11090 8250 11110 8320
rect 11180 8250 11200 8320
rect 11270 8250 11290 8320
rect 11360 8250 11380 8320
rect 11450 8250 11470 8320
rect 11540 8250 11560 8320
rect 11630 8250 11650 8320
rect 11720 8250 11740 8320
rect 11810 8250 11830 8320
rect 11900 8250 11920 8320
rect 11990 8250 12010 8320
rect 12080 8250 12100 8320
rect 12170 8250 12190 8320
rect 12260 8250 12280 8320
rect 12350 8250 12370 8320
rect 12440 8250 12460 8320
rect 12530 8250 12550 8320
rect 12620 8250 12640 8320
rect 12710 8250 12730 8320
rect 12800 8250 12820 8320
rect 12890 8250 12910 8320
rect 12980 8250 13000 8320
rect 13070 8250 13090 8320
rect 13160 8250 13180 8320
rect 13250 8250 13270 8320
rect 13340 8250 13360 8320
rect 13430 8250 13450 8320
rect 13520 8250 13540 8320
rect 13610 8250 13670 8320
rect 13740 8250 13760 8320
rect 13830 8250 13850 8320
rect 13920 8250 13940 8320
rect 14010 8250 14030 8320
rect 14100 8250 14120 8320
rect 14190 8250 14210 8320
rect 14280 8250 14300 8320
rect 14370 8250 14390 8320
rect 14460 8250 14480 8320
rect 14550 8250 14570 8320
rect 14640 8250 14660 8320
rect 14730 8250 14750 8320
rect 14820 8250 14840 8320
rect 14910 8250 14930 8320
rect 15000 8250 15020 8320
rect 15090 8250 15110 8320
rect 15180 8250 15200 8320
rect 15270 8250 15290 8320
rect 15360 8250 15380 8320
rect 15450 8250 15470 8320
rect 15540 8250 15560 8320
rect 15630 8250 15650 8320
rect 15720 8250 15740 8320
rect 15810 8250 15830 8320
rect 15900 8250 15920 8320
rect 15990 8250 16010 8320
rect 16080 8250 16100 8320
rect 16170 8250 16190 8320
rect 16260 8250 16280 8320
rect 16350 8250 16370 8320
rect 16440 8250 16460 8320
rect 16530 8250 16550 8320
rect 16620 8250 16680 8320
rect 16750 8250 16770 8320
rect 16840 8250 16860 8320
rect 16930 8250 16950 8320
rect 17020 8250 17040 8320
rect 17110 8250 17130 8320
rect 17200 8250 17220 8320
rect 17290 8250 17310 8320
rect 17380 8250 17400 8320
rect 17470 8250 17490 8320
rect 17560 8250 17580 8320
rect 17650 8250 17670 8320
rect 17740 8250 17760 8320
rect 17830 8250 17850 8320
rect 17920 8250 17940 8320
rect 18010 8250 18030 8320
rect 18100 8250 18120 8320
rect 18190 8250 18210 8320
rect 18280 8250 18300 8320
rect 18370 8250 18390 8320
rect 18460 8250 18480 8320
rect 18550 8250 18570 8320
rect 18640 8250 18660 8320
rect 18730 8250 18750 8320
rect 18820 8250 18840 8320
rect 18910 8250 18930 8320
rect 19000 8250 19020 8320
rect 19090 8250 19110 8320
rect 19180 8250 19200 8320
rect 19270 8250 19290 8320
rect 19360 8250 19380 8320
rect 19450 8250 19470 8320
rect 19540 8250 19560 8320
rect 19630 8250 19920 8320
rect 7610 8190 19920 8250
rect 7020 7910 7340 7930
rect 7020 7840 7040 7910
rect 7110 7840 7140 7910
rect 7210 7840 7240 7910
rect 7310 7840 7340 7910
rect 7020 7820 7340 7840
rect 7020 7750 7040 7820
rect 7110 7750 7140 7820
rect 7210 7750 7240 7820
rect 7310 7750 7340 7820
rect 1540 6850 3140 6900
rect 1540 6780 1570 6850
rect 1640 6780 1680 6850
rect 1750 6780 1790 6850
rect 1860 6780 1900 6850
rect 1970 6780 2010 6850
rect 2080 6780 2120 6850
rect 2190 6780 2230 6850
rect 2300 6780 2340 6850
rect 2410 6780 2450 6850
rect 2520 6780 2560 6850
rect 2630 6780 2670 6850
rect 2740 6780 2780 6850
rect 2850 6780 2890 6850
rect 2960 6780 3000 6850
rect 3070 6780 3140 6850
rect 1540 6740 3140 6780
rect 1540 6670 1570 6740
rect 1640 6670 1680 6740
rect 1750 6670 1790 6740
rect 1860 6670 1900 6740
rect 1970 6670 2010 6740
rect 2080 6670 2120 6740
rect 2190 6670 2230 6740
rect 2300 6670 2340 6740
rect 2410 6670 2450 6740
rect 2520 6670 2560 6740
rect 2630 6670 2670 6740
rect 2740 6670 2780 6740
rect 2850 6670 2890 6740
rect 2960 6670 3000 6740
rect 3070 6670 3140 6740
rect 1540 6640 3140 6670
rect 7020 4610 7340 7750
rect 7560 7910 7880 7930
rect 7560 7840 7590 7910
rect 7660 7840 7690 7910
rect 7760 7840 7790 7910
rect 7860 7840 7880 7910
rect 7560 7820 7880 7840
rect 7560 7750 7590 7820
rect 7660 7750 7690 7820
rect 7760 7750 7790 7820
rect 7860 7750 7880 7820
rect 7400 5390 7490 5410
rect 7400 5320 7410 5390
rect 7480 5320 7490 5390
rect 7400 5280 7490 5320
rect 7400 5210 7410 5280
rect 7480 5210 7490 5280
rect 7400 5170 7490 5210
rect 7400 5100 7410 5170
rect 7480 5100 7490 5170
rect 7400 5060 7490 5100
rect 7400 4990 7410 5060
rect 7480 4990 7490 5060
rect 7400 4950 7490 4990
rect 7400 4880 7410 4950
rect 7480 4880 7490 4950
rect 7400 4860 7490 4880
rect 7560 4760 7880 7750
rect 28700 7820 36100 7910
rect 28700 7750 35790 7820
rect 35860 7750 35880 7820
rect 35950 7750 35970 7820
rect 36040 7750 36100 7820
rect 28700 7730 36100 7750
rect 28700 7660 35790 7730
rect 35860 7660 35880 7730
rect 35950 7660 35970 7730
rect 36040 7660 36100 7730
rect 28700 7640 36100 7660
rect 28700 7570 35790 7640
rect 35860 7570 35880 7640
rect 35950 7570 35970 7640
rect 36040 7570 36100 7640
rect 28700 7550 36100 7570
rect 28700 7480 35790 7550
rect 35860 7480 35880 7550
rect 35950 7480 35970 7550
rect 36040 7480 36100 7550
rect 28700 7460 36100 7480
rect 28700 7390 35790 7460
rect 35860 7390 35880 7460
rect 35950 7390 35970 7460
rect 36040 7390 36100 7460
rect 28700 7370 36100 7390
rect 28700 7300 35790 7370
rect 35860 7300 35880 7370
rect 35950 7300 35970 7370
rect 36040 7300 36100 7370
rect 28700 7280 36100 7300
rect 21060 7210 21540 7260
rect 21060 7140 21090 7210
rect 21160 7140 21200 7210
rect 21270 7140 21310 7210
rect 21380 7140 21420 7210
rect 21490 7140 21540 7210
rect 21060 7100 21540 7140
rect 21060 7030 21090 7100
rect 21160 7030 21200 7100
rect 21270 7030 21310 7100
rect 21380 7030 21420 7100
rect 21490 7030 21540 7100
rect 21060 7000 21540 7030
rect 23460 7210 23940 7260
rect 23460 7140 23490 7210
rect 23560 7140 23600 7210
rect 23670 7140 23710 7210
rect 23780 7140 23820 7210
rect 23890 7140 23940 7210
rect 23460 7100 23940 7140
rect 23460 7030 23490 7100
rect 23560 7030 23600 7100
rect 23670 7030 23710 7100
rect 23780 7030 23820 7100
rect 23890 7030 23940 7100
rect 23460 7000 23940 7030
rect 28700 7210 35790 7280
rect 35860 7210 35880 7280
rect 35950 7210 35970 7280
rect 36040 7210 36100 7280
rect 28700 7150 36100 7210
rect 28700 7080 35790 7150
rect 35860 7080 35880 7150
rect 35950 7080 35970 7150
rect 36040 7080 36100 7150
rect 28700 7060 36100 7080
rect 28700 6990 35790 7060
rect 35860 6990 35880 7060
rect 35950 6990 35970 7060
rect 36040 6990 36100 7060
rect 28700 6970 36100 6990
rect 11760 6880 13360 6930
rect 11760 6810 11790 6880
rect 11860 6810 11900 6880
rect 11970 6810 12010 6880
rect 12080 6810 12120 6880
rect 12190 6810 12230 6880
rect 12300 6810 12340 6880
rect 12410 6810 12450 6880
rect 12520 6810 12560 6880
rect 12630 6810 12670 6880
rect 12740 6810 12780 6880
rect 12850 6810 12890 6880
rect 12960 6810 13000 6880
rect 13070 6810 13110 6880
rect 13180 6810 13220 6880
rect 13290 6810 13360 6880
rect 11760 6770 13360 6810
rect 11760 6700 11790 6770
rect 11860 6700 11900 6770
rect 11970 6700 12010 6770
rect 12080 6700 12120 6770
rect 12190 6700 12230 6770
rect 12300 6700 12340 6770
rect 12410 6700 12450 6770
rect 12520 6700 12560 6770
rect 12630 6700 12670 6770
rect 12740 6700 12780 6770
rect 12850 6700 12890 6770
rect 12960 6700 13000 6770
rect 13070 6700 13110 6770
rect 13180 6700 13220 6770
rect 13290 6700 13360 6770
rect 11760 6670 13360 6700
rect 28700 6900 35790 6970
rect 35860 6900 35880 6970
rect 35950 6900 35970 6970
rect 36040 6900 36100 6970
rect 28700 6880 36100 6900
rect 28700 6810 35790 6880
rect 35860 6810 35880 6880
rect 35950 6810 35970 6880
rect 36040 6810 36100 6880
rect 28700 6790 36100 6810
rect 28700 6720 35790 6790
rect 35860 6720 35880 6790
rect 35950 6720 35970 6790
rect 36040 6720 36100 6790
rect 28700 6700 36100 6720
rect 28700 6630 35790 6700
rect 35860 6630 35880 6700
rect 35950 6630 35970 6700
rect 36040 6630 36100 6700
rect 28700 6610 36100 6630
rect 28700 6540 35790 6610
rect 35860 6540 35880 6610
rect 35950 6540 35970 6610
rect 36040 6540 36100 6610
rect 28700 6520 36100 6540
rect 28700 6450 35790 6520
rect 35860 6450 35880 6520
rect 35950 6450 35970 6520
rect 36040 6450 36100 6520
rect 28700 6430 36100 6450
rect 28700 6360 35790 6430
rect 35860 6360 35880 6430
rect 35950 6360 35970 6430
rect 36040 6360 36100 6430
rect 28700 6340 36100 6360
rect 28320 6300 28540 6320
rect 28320 6230 28340 6300
rect 28410 6230 28450 6300
rect 28520 6230 28540 6300
rect 28320 6170 28540 6230
rect 28320 6100 28340 6170
rect 28410 6100 28450 6170
rect 28520 6100 28540 6170
rect 28320 6040 28540 6100
rect 28320 5970 28340 6040
rect 28410 5970 28450 6040
rect 28520 5970 28540 6040
rect 28320 5950 28540 5970
rect 28700 6270 35790 6340
rect 35860 6270 35880 6340
rect 35950 6270 35970 6340
rect 36040 6270 36100 6340
rect 28700 6250 36100 6270
rect 28700 6180 35790 6250
rect 35860 6180 35880 6250
rect 35950 6180 35970 6250
rect 36040 6180 36100 6250
rect 28700 6160 36100 6180
rect 28700 6090 35790 6160
rect 35860 6090 35880 6160
rect 35950 6090 35970 6160
rect 36040 6090 36100 6160
rect 28700 6070 36100 6090
rect 28700 6000 35790 6070
rect 35860 6000 35880 6070
rect 35950 6000 35970 6070
rect 36040 6000 36100 6070
rect 28700 5980 36100 6000
rect 7560 4700 7590 4760
rect 7650 4700 7690 4760
rect 7750 4700 7790 4760
rect 7850 4700 7880 4760
rect 7560 4670 7880 4700
rect 28700 5910 35790 5980
rect 35860 5910 35880 5980
rect 35950 5910 35970 5980
rect 36040 5910 36100 5980
rect 28700 5890 36100 5910
rect 28700 5820 35790 5890
rect 35860 5820 35880 5890
rect 35950 5820 35970 5890
rect 36040 5820 36100 5890
rect 28700 5800 36100 5820
rect 28700 5730 35790 5800
rect 35860 5730 35880 5800
rect 35950 5730 35970 5800
rect 36040 5730 36100 5800
rect 28700 5710 36100 5730
rect 28700 5640 35790 5710
rect 35860 5640 35880 5710
rect 35950 5640 35970 5710
rect 36040 5640 36100 5710
rect 28700 5620 36100 5640
rect 28700 5550 35790 5620
rect 35860 5550 35880 5620
rect 35950 5550 35970 5620
rect 36040 5550 36100 5620
rect 28700 5530 36100 5550
rect 28700 5460 35790 5530
rect 35860 5460 35880 5530
rect 35950 5460 35970 5530
rect 36040 5460 36100 5530
rect 28700 5440 36100 5460
rect 28700 5370 35790 5440
rect 35860 5370 35880 5440
rect 35950 5370 35970 5440
rect 36040 5370 36100 5440
rect 28700 5350 36100 5370
rect 28700 5280 35790 5350
rect 35860 5280 35880 5350
rect 35950 5280 35970 5350
rect 36040 5280 36100 5350
rect 28700 5260 36100 5280
rect 28700 5190 35790 5260
rect 35860 5190 35880 5260
rect 35950 5190 35970 5260
rect 36040 5190 36100 5260
rect 28700 5170 36100 5190
rect 28700 5100 35790 5170
rect 35860 5100 35880 5170
rect 35950 5100 35970 5170
rect 36040 5100 36100 5170
rect 28700 5080 36100 5100
rect 28700 5010 35790 5080
rect 35860 5010 35880 5080
rect 35950 5010 35970 5080
rect 36040 5010 36100 5080
rect 28700 4990 36100 5010
rect 28700 4920 35790 4990
rect 35860 4920 35880 4990
rect 35950 4920 35970 4990
rect 36040 4920 36100 4990
rect 28700 4900 36100 4920
rect 28700 4830 35790 4900
rect 35860 4830 35880 4900
rect 35950 4830 35970 4900
rect 36040 4830 36100 4900
rect 28700 4810 36100 4830
rect 28700 4740 35790 4810
rect 35860 4740 35880 4810
rect 35950 4740 35970 4810
rect 36040 4740 36100 4810
rect 28700 4720 36100 4740
rect 28700 4650 35790 4720
rect 35860 4650 35880 4720
rect 35950 4650 35970 4720
rect 36040 4650 36100 4720
rect 28700 4630 36100 4650
rect -880 4580 6790 4610
rect -880 4510 -840 4580
rect -770 4510 -710 4580
rect -640 4520 6700 4580
rect 6760 4520 6790 4580
rect -640 4510 6790 4520
rect -880 4470 6790 4510
rect -880 4400 -840 4470
rect -770 4400 -710 4470
rect -640 4460 6790 4470
rect -640 4400 6700 4460
rect 6760 4400 6790 4460
rect -880 4360 6790 4400
rect -880 4290 -840 4360
rect -770 4290 -710 4360
rect -640 4340 6790 4360
rect -640 4290 6700 4340
rect -880 4280 6700 4290
rect 6760 4280 6790 4340
rect -880 4250 6790 4280
rect -880 4180 -840 4250
rect -770 4180 -710 4250
rect -640 4220 6790 4250
rect -640 4180 6700 4220
rect -880 4160 6700 4180
rect 6760 4160 6790 4220
rect -880 4130 6790 4160
rect 7020 4580 15660 4610
rect 7020 4510 15420 4580
rect 15490 4510 15550 4580
rect 15620 4510 15660 4580
rect 7020 4470 15660 4510
rect 7020 4400 15420 4470
rect 15490 4400 15550 4470
rect 15620 4400 15660 4470
rect 7020 4360 15660 4400
rect 7020 4290 15420 4360
rect 15490 4290 15550 4360
rect 15620 4290 15660 4360
rect 7020 4250 15660 4290
rect 7020 4180 15420 4250
rect 15490 4180 15550 4250
rect 15620 4180 15660 4250
rect 7020 4130 15660 4180
rect 28700 4560 35790 4630
rect 35860 4560 35880 4630
rect 35950 4560 35970 4630
rect 36040 4560 36100 4630
rect 28700 4540 36100 4560
rect 28700 4470 35790 4540
rect 35860 4470 35880 4540
rect 35950 4470 35970 4540
rect 36040 4470 36100 4540
rect 28700 4450 36100 4470
rect 28700 4380 35790 4450
rect 35860 4380 35880 4450
rect 35950 4380 35970 4450
rect 36040 4380 36100 4450
rect 28700 4360 36100 4380
rect 28700 4290 35790 4360
rect 35860 4290 35880 4360
rect 35950 4290 35970 4360
rect 36040 4290 36100 4360
rect 28700 4270 36100 4290
rect 28700 4200 35790 4270
rect 35860 4200 35880 4270
rect 35950 4200 35970 4270
rect 36040 4200 36100 4270
rect 28700 4140 36100 4200
rect 7020 3240 7340 4130
rect 28700 4070 35790 4140
rect 35860 4070 35880 4140
rect 35950 4070 35970 4140
rect 36040 4070 36100 4140
rect 28700 4050 36100 4070
rect 28700 3980 35790 4050
rect 35860 3980 35880 4050
rect 35950 3980 35970 4050
rect 36040 3980 36100 4050
rect 28700 3960 36100 3980
rect 28700 3890 35790 3960
rect 35860 3890 35880 3960
rect 35950 3890 35970 3960
rect 36040 3890 36100 3960
rect 28700 3870 36100 3890
rect 28700 3800 35790 3870
rect 35860 3800 35880 3870
rect 35950 3800 35970 3870
rect 36040 3800 36100 3870
rect 28700 3780 36100 3800
rect 28700 3710 35790 3780
rect 35860 3710 35880 3780
rect 35950 3710 35970 3780
rect 36040 3710 36100 3780
rect 28700 3690 36100 3710
rect 28700 3620 35790 3690
rect 35860 3620 35880 3690
rect 35950 3620 35970 3690
rect 36040 3620 36100 3690
rect 28700 3600 36100 3620
rect 28700 3530 35790 3600
rect 35860 3530 35880 3600
rect 35950 3530 35970 3600
rect 36040 3530 36100 3600
rect 28700 3510 36100 3530
rect 28700 3440 35790 3510
rect 35860 3440 35880 3510
rect 35950 3440 35970 3510
rect 36040 3440 36100 3510
rect 28700 3420 36100 3440
rect 7020 3180 7050 3240
rect 7110 3180 7150 3240
rect 7210 3180 7250 3240
rect 7310 3180 7340 3240
rect 7020 3140 7340 3180
rect 7020 3080 7050 3140
rect 7110 3080 7150 3140
rect 7210 3080 7250 3140
rect 7310 3080 7340 3140
rect 7020 3040 7340 3080
rect 22300 3360 22630 3380
rect 22300 3290 22320 3360
rect 22390 3290 22430 3360
rect 22500 3290 22540 3360
rect 22610 3290 22630 3360
rect 22300 3250 22630 3290
rect 22300 3180 22320 3250
rect 22390 3180 22430 3250
rect 22500 3180 22540 3250
rect 22610 3180 22630 3250
rect 22300 3140 22630 3180
rect 22300 3070 22320 3140
rect 22390 3070 22430 3140
rect 22500 3070 22540 3140
rect 22610 3070 22630 3140
rect 22300 3050 22630 3070
rect 28700 3350 35790 3420
rect 35860 3350 35880 3420
rect 35950 3350 35970 3420
rect 36040 3350 36100 3420
rect 28700 3330 36100 3350
rect 28700 3260 35790 3330
rect 35860 3260 35880 3330
rect 35950 3260 35970 3330
rect 36040 3260 36100 3330
rect 28700 3240 36100 3260
rect 28700 3170 35790 3240
rect 35860 3170 35880 3240
rect 35950 3170 35970 3240
rect 36040 3170 36100 3240
rect 28700 3150 36100 3170
rect 28700 3080 35790 3150
rect 35860 3080 35880 3150
rect 35950 3080 35970 3150
rect 36040 3080 36100 3150
rect 28700 3060 36100 3080
rect 7020 2980 7050 3040
rect 7110 2980 7150 3040
rect 7210 2980 7250 3040
rect 7310 2980 7340 3040
rect 7020 2960 7340 2980
rect 28700 2990 35790 3060
rect 35860 2990 35880 3060
rect 35950 2990 35970 3060
rect 36040 2990 36100 3060
rect 28700 2970 36100 2990
rect 4740 2890 6750 2920
rect 4740 2830 4770 2890
rect 4830 2830 4870 2890
rect 4930 2830 4970 2890
rect 5030 2830 6750 2890
rect 4740 2790 6750 2830
rect 4740 2730 4770 2790
rect 4830 2730 4870 2790
rect 4930 2730 4970 2790
rect 5030 2730 6750 2790
rect 4740 2690 6750 2730
rect 4740 2630 4770 2690
rect 4830 2630 4870 2690
rect 4930 2630 4970 2690
rect 5030 2630 6750 2690
rect 4740 2610 6750 2630
rect 6440 -100 6750 2610
rect -330 -140 6750 -100
rect -330 -210 -300 -140
rect -230 -210 -190 -140
rect -120 -210 -80 -140
rect -10 -210 30 -140
rect 100 -210 6750 -140
rect -330 -270 6750 -210
rect -330 -340 -300 -270
rect -230 -340 -190 -270
rect -120 -340 -80 -270
rect -10 -340 30 -270
rect 100 -340 6750 -270
rect -330 -380 6750 -340
rect 1080 -790 2680 -760
rect 1080 -860 1150 -790
rect 1220 -860 1260 -790
rect 1330 -860 1370 -790
rect 1440 -860 1480 -790
rect 1550 -860 1590 -790
rect 1660 -860 1700 -790
rect 1770 -860 1810 -790
rect 1880 -860 1920 -790
rect 1990 -860 2030 -790
rect 2100 -860 2140 -790
rect 2210 -860 2250 -790
rect 2320 -860 2360 -790
rect 2430 -860 2470 -790
rect 2540 -860 2580 -790
rect 2650 -860 2680 -790
rect 1080 -900 2680 -860
rect 1080 -970 1150 -900
rect 1220 -970 1260 -900
rect 1330 -970 1370 -900
rect 1440 -970 1480 -900
rect 1550 -970 1590 -900
rect 1660 -970 1700 -900
rect 1770 -970 1810 -900
rect 1880 -970 1920 -900
rect 1990 -970 2030 -900
rect 2100 -970 2140 -900
rect 2210 -970 2250 -900
rect 2320 -970 2360 -900
rect 2430 -970 2470 -900
rect 2540 -970 2580 -900
rect 2650 -970 2680 -900
rect 1080 -1020 2680 -970
rect 1540 -2780 3140 -2730
rect 1540 -2850 1570 -2780
rect 1640 -2850 1680 -2780
rect 1750 -2850 1790 -2780
rect 1860 -2850 1900 -2780
rect 1970 -2850 2010 -2780
rect 2080 -2850 2120 -2780
rect 2190 -2850 2230 -2780
rect 2300 -2850 2340 -2780
rect 2410 -2850 2450 -2780
rect 2520 -2850 2560 -2780
rect 2630 -2850 2670 -2780
rect 2740 -2850 2780 -2780
rect 2850 -2850 2890 -2780
rect 2960 -2850 3000 -2780
rect 3070 -2850 3140 -2780
rect 1540 -2890 3140 -2850
rect 1540 -2960 1570 -2890
rect 1640 -2960 1680 -2890
rect 1750 -2960 1790 -2890
rect 1860 -2960 1900 -2890
rect 1970 -2960 2010 -2890
rect 2080 -2960 2120 -2890
rect 2190 -2960 2230 -2890
rect 2300 -2960 2340 -2890
rect 2410 -2960 2450 -2890
rect 2520 -2960 2560 -2890
rect 2630 -2960 2670 -2890
rect 2740 -2960 2780 -2890
rect 2850 -2960 2890 -2890
rect 2960 -2960 3000 -2890
rect 3070 -2960 3140 -2890
rect 1540 -2990 3140 -2960
rect 6440 -3700 6750 -380
rect -2220 -3970 6750 -3700
rect -2220 -4470 -1940 -3970
rect -2220 -4540 -2200 -4470
rect -2130 -4540 -2090 -4470
rect -2020 -4540 -1940 -4470
rect -2220 -4580 -1940 -4540
rect -2220 -4650 -2200 -4580
rect -2130 -4650 -2090 -4580
rect -2020 -4650 -1940 -4580
rect -2220 -4690 -1940 -4650
rect -2220 -4760 -2200 -4690
rect -2130 -4760 -2090 -4690
rect -2020 -4760 -1940 -4690
rect -2220 -4800 -1940 -4760
rect -2220 -4870 -2200 -4800
rect -2130 -4870 -2090 -4800
rect -2020 -4870 -1940 -4800
rect -2220 -4900 -1940 -4870
rect -1860 -4230 150 -4050
rect -1860 -4300 -160 -4230
rect -90 -4300 -70 -4230
rect 0 -4300 20 -4230
rect 90 -4300 150 -4230
rect -1860 -4320 150 -4300
rect -1860 -4390 -160 -4320
rect -90 -4390 -70 -4320
rect 0 -4390 20 -4320
rect 90 -4390 150 -4320
rect -1860 -4410 150 -4390
rect -1860 -4480 -160 -4410
rect -90 -4480 -70 -4410
rect 0 -4480 20 -4410
rect 90 -4480 150 -4410
rect -1860 -4500 150 -4480
rect -1860 -4570 -160 -4500
rect -90 -4570 -70 -4500
rect 0 -4570 20 -4500
rect 90 -4570 150 -4500
rect -1860 -4590 150 -4570
rect -1860 -4660 -160 -4590
rect -90 -4660 -70 -4590
rect 0 -4660 20 -4590
rect 90 -4660 150 -4590
rect -1860 -4680 150 -4660
rect -1860 -4750 -160 -4680
rect -90 -4750 -70 -4680
rect 0 -4750 20 -4680
rect 90 -4750 150 -4680
rect -1860 -4770 150 -4750
rect -1860 -4840 -160 -4770
rect -90 -4840 -70 -4770
rect 0 -4840 20 -4770
rect 90 -4840 150 -4770
rect -1860 -4860 150 -4840
rect -1860 -4930 -160 -4860
rect -90 -4930 -70 -4860
rect 0 -4930 20 -4860
rect 90 -4930 150 -4860
rect -1860 -4950 150 -4930
rect -1860 -5020 -160 -4950
rect -90 -5020 -70 -4950
rect 0 -5020 20 -4950
rect 90 -5020 150 -4950
rect -1860 -5040 150 -5020
rect -1860 -5110 -160 -5040
rect -90 -5110 -70 -5040
rect 0 -5110 20 -5040
rect 90 -5110 150 -5040
rect -1860 -5130 150 -5110
rect -1860 -5200 -160 -5130
rect -90 -5200 -70 -5130
rect 0 -5200 20 -5130
rect 90 -5200 150 -5130
rect -1860 -5220 150 -5200
rect -2160 -5240 -1940 -5220
rect -2160 -5310 -2140 -5240
rect -2070 -5310 -2030 -5240
rect -1960 -5310 -1940 -5240
rect -2160 -5350 -1940 -5310
rect -2160 -5420 -2140 -5350
rect -2070 -5420 -2030 -5350
rect -1960 -5420 -1940 -5350
rect -2160 -5460 -1940 -5420
rect -2160 -5530 -2140 -5460
rect -2070 -5530 -2030 -5460
rect -1960 -5530 -1940 -5460
rect -2160 -5570 -1940 -5530
rect -2160 -5640 -2140 -5570
rect -2070 -5640 -2030 -5570
rect -1960 -5640 -1940 -5570
rect -2160 -5660 -1940 -5640
rect -1860 -5290 -160 -5220
rect -90 -5290 -70 -5220
rect 0 -5290 20 -5220
rect 90 -5290 150 -5220
rect -1860 -5310 150 -5290
rect -1860 -5380 -160 -5310
rect -90 -5380 -70 -5310
rect 0 -5380 20 -5310
rect 90 -5380 150 -5310
rect -1860 -5400 150 -5380
rect -1860 -5470 -160 -5400
rect -90 -5470 -70 -5400
rect 0 -5470 20 -5400
rect 90 -5470 150 -5400
rect -1860 -5660 150 -5470
rect -880 -6500 -600 -6470
rect -880 -6570 -840 -6500
rect -770 -6570 -710 -6500
rect -640 -6570 -600 -6500
rect -880 -6610 -600 -6570
rect -880 -6680 -840 -6610
rect -770 -6680 -710 -6610
rect -640 -6640 -600 -6610
rect -180 -6640 150 -5660
rect 6440 -6420 6750 -3970
rect 8180 2890 10160 2920
rect 8180 2830 9870 2890
rect 9930 2830 9970 2890
rect 10030 2830 10070 2890
rect 10130 2830 10160 2890
rect 8180 2790 10160 2830
rect 8180 2730 9870 2790
rect 9930 2730 9970 2790
rect 10030 2730 10070 2790
rect 10130 2730 10160 2790
rect 8180 2690 10160 2730
rect 8180 2630 9870 2690
rect 9930 2630 9970 2690
rect 10030 2630 10070 2690
rect 10130 2630 10160 2690
rect 28700 2900 35790 2970
rect 35860 2900 35880 2970
rect 35950 2900 35970 2970
rect 36040 2900 36100 2970
rect 28700 2880 36100 2900
rect 28700 2810 35790 2880
rect 35860 2810 35880 2880
rect 35950 2810 35970 2880
rect 36040 2810 36100 2880
rect 28700 2790 36100 2810
rect 28700 2720 35790 2790
rect 35860 2720 35880 2790
rect 35950 2720 35970 2790
rect 36040 2720 36100 2790
rect 28700 2700 36100 2720
rect 28700 2630 35790 2700
rect 35860 2630 35880 2700
rect 35950 2630 35970 2700
rect 36040 2630 36100 2700
rect 8180 2610 10160 2630
rect 8180 -100 8490 2610
rect 20020 2600 20500 2630
rect 20020 2530 20070 2600
rect 20140 2530 20180 2600
rect 20250 2530 20290 2600
rect 20360 2530 20400 2600
rect 20470 2530 20500 2600
rect 20020 2490 20500 2530
rect 20020 2420 20070 2490
rect 20140 2420 20180 2490
rect 20250 2420 20290 2490
rect 20360 2420 20400 2490
rect 20470 2420 20500 2490
rect 20020 2370 20500 2420
rect 24500 2600 24980 2630
rect 24500 2530 24550 2600
rect 24620 2530 24660 2600
rect 24730 2530 24770 2600
rect 24840 2530 24880 2600
rect 24950 2530 24980 2600
rect 24500 2490 24980 2530
rect 24500 2420 24550 2490
rect 24620 2420 24660 2490
rect 24730 2420 24770 2490
rect 24840 2420 24880 2490
rect 24950 2420 24980 2490
rect 24500 2370 24980 2420
rect 28700 2610 36100 2630
rect 28700 2540 35790 2610
rect 35860 2540 35880 2610
rect 35950 2540 35970 2610
rect 36040 2540 36100 2610
rect 28700 2520 36100 2540
rect 28700 2450 35790 2520
rect 35860 2450 35880 2520
rect 35950 2450 35970 2520
rect 36040 2450 36100 2520
rect 28700 2430 36100 2450
rect 28700 2360 35790 2430
rect 35860 2360 35880 2430
rect 35950 2360 35970 2430
rect 36040 2360 36100 2430
rect 28700 2340 36100 2360
rect 28700 2270 35790 2340
rect 35860 2270 35880 2340
rect 35950 2270 35970 2340
rect 36040 2270 36100 2340
rect 28700 2250 36100 2270
rect 28700 2180 35790 2250
rect 35860 2180 35880 2250
rect 35950 2180 35970 2250
rect 36040 2180 36100 2250
rect 28700 2160 36100 2180
rect 28700 2090 35790 2160
rect 35860 2090 35880 2160
rect 35950 2090 35970 2160
rect 36040 2090 36100 2160
rect 28700 2070 36100 2090
rect 28700 2000 35790 2070
rect 35860 2000 35880 2070
rect 35950 2000 35970 2070
rect 36040 2000 36100 2070
rect 28700 1980 36100 2000
rect 28700 1910 35790 1980
rect 35860 1910 35880 1980
rect 35950 1910 35970 1980
rect 36040 1910 36100 1980
rect 28700 1890 36100 1910
rect 28700 1820 35790 1890
rect 35860 1820 35880 1890
rect 35950 1820 35970 1890
rect 36040 1820 36100 1890
rect 28700 1800 36100 1820
rect 28700 1730 35790 1800
rect 35860 1730 35880 1800
rect 35950 1730 35970 1800
rect 36040 1730 36100 1800
rect 28700 1710 36100 1730
rect 28700 1640 35790 1710
rect 35860 1640 35880 1710
rect 35950 1640 35970 1710
rect 36040 1640 36100 1710
rect 28700 1620 36100 1640
rect 28700 1550 35790 1620
rect 35860 1550 35880 1620
rect 35950 1550 35970 1620
rect 36040 1550 36100 1620
rect 28700 1530 36100 1550
rect 28700 1460 35790 1530
rect 35860 1460 35880 1530
rect 35950 1460 35970 1530
rect 36040 1460 36100 1530
rect 28700 1440 36100 1460
rect 28700 1370 35790 1440
rect 35860 1370 35880 1440
rect 35950 1370 35970 1440
rect 36040 1370 36100 1440
rect 28700 1350 36100 1370
rect 28700 1280 35790 1350
rect 35860 1280 35880 1350
rect 35950 1280 35970 1350
rect 36040 1280 36100 1350
rect 28700 1260 36100 1280
rect 28700 1190 35790 1260
rect 35860 1190 35880 1260
rect 35950 1190 35970 1260
rect 36040 1190 36100 1260
rect 14590 1160 14900 1180
rect 14590 1090 14600 1160
rect 14670 1090 14700 1160
rect 14770 1090 14810 1160
rect 14880 1090 14900 1160
rect 28700 1150 36100 1190
rect 14590 1050 14900 1090
rect 14590 980 14600 1050
rect 14670 980 14700 1050
rect 14770 980 14810 1050
rect 14880 980 14900 1050
rect 14590 940 14900 980
rect 14590 870 14600 940
rect 14670 870 14700 940
rect 14770 870 14810 940
rect 14880 870 14900 940
rect 14590 850 14900 870
rect 21060 920 21540 970
rect 21060 850 21090 920
rect 21160 850 21200 920
rect 21270 850 21310 920
rect 21380 850 21420 920
rect 21490 850 21540 920
rect 21060 810 21540 850
rect 21060 740 21090 810
rect 21160 740 21200 810
rect 21270 740 21310 810
rect 21380 740 21420 810
rect 21490 740 21540 810
rect 21060 710 21540 740
rect 23460 920 23940 970
rect 23460 850 23490 920
rect 23560 850 23600 920
rect 23670 850 23710 920
rect 23780 850 23820 920
rect 23890 850 23940 920
rect 23460 810 23940 850
rect 23460 740 23490 810
rect 23560 740 23600 810
rect 23670 740 23710 810
rect 23780 740 23820 810
rect 23890 740 23940 810
rect 23460 710 23940 740
rect 28700 220 36100 310
rect 28700 150 35790 220
rect 35860 150 35880 220
rect 35950 150 35970 220
rect 36040 150 36100 220
rect 28700 130 36100 150
rect 28700 60 35790 130
rect 35860 60 35880 130
rect 35950 60 35970 130
rect 36040 60 36100 130
rect 28700 40 36100 60
rect 28320 0 28540 20
rect 28320 -70 28340 0
rect 28410 -70 28450 0
rect 28520 -70 28540 0
rect 8180 -140 15110 -100
rect 8180 -210 14660 -140
rect 14730 -210 14770 -140
rect 14840 -210 14880 -140
rect 14950 -210 14990 -140
rect 15060 -210 15110 -140
rect 8180 -270 15110 -210
rect 8180 -340 14660 -270
rect 14730 -340 14770 -270
rect 14840 -340 14880 -270
rect 14950 -340 14990 -270
rect 15060 -340 15110 -270
rect 8180 -380 15110 -340
rect 28320 -130 28540 -70
rect 28320 -200 28340 -130
rect 28410 -200 28450 -130
rect 28520 -200 28540 -130
rect 28320 -260 28540 -200
rect 28320 -330 28340 -260
rect 28410 -330 28450 -260
rect 28520 -330 28540 -260
rect 28320 -350 28540 -330
rect 28700 -30 35790 40
rect 35860 -30 35880 40
rect 35950 -30 35970 40
rect 36040 -30 36100 40
rect 28700 -50 36100 -30
rect 28700 -120 35790 -50
rect 35860 -120 35880 -50
rect 35950 -120 35970 -50
rect 36040 -120 36100 -50
rect 28700 -140 36100 -120
rect 28700 -210 35790 -140
rect 35860 -210 35880 -140
rect 35950 -210 35970 -140
rect 36040 -210 36100 -140
rect 28700 -230 36100 -210
rect 28700 -300 35790 -230
rect 35860 -300 35880 -230
rect 35950 -300 35970 -230
rect 36040 -300 36100 -230
rect 28700 -320 36100 -300
rect 7290 -4560 7620 -4540
rect 7290 -4630 7310 -4560
rect 7380 -4630 7420 -4560
rect 7490 -4630 7530 -4560
rect 7600 -4630 7620 -4560
rect 7290 -4670 7620 -4630
rect 7290 -4740 7310 -4670
rect 7380 -4740 7420 -4670
rect 7490 -4740 7530 -4670
rect 7600 -4740 7620 -4670
rect 7290 -4780 7620 -4740
rect 7290 -4850 7310 -4780
rect 7380 -4850 7420 -4780
rect 7490 -4850 7530 -4780
rect 7600 -4850 7620 -4780
rect 7290 -4870 7620 -4850
rect 8180 -6150 8490 -380
rect 28700 -390 35790 -320
rect 35860 -390 35880 -320
rect 35950 -390 35970 -320
rect 36040 -390 36100 -320
rect 28700 -450 36100 -390
rect 28700 -520 35790 -450
rect 35860 -520 35880 -450
rect 35950 -520 35970 -450
rect 36040 -520 36100 -450
rect 28700 -540 36100 -520
rect 28700 -610 35790 -540
rect 35860 -610 35880 -540
rect 35950 -610 35970 -540
rect 36040 -610 36100 -540
rect 28700 -630 36100 -610
rect 28700 -700 35790 -630
rect 35860 -700 35880 -630
rect 35950 -700 35970 -630
rect 36040 -700 36100 -630
rect 28700 -720 36100 -700
rect 12220 -790 13820 -760
rect 12220 -860 12250 -790
rect 12320 -860 12360 -790
rect 12430 -860 12470 -790
rect 12540 -860 12580 -790
rect 12650 -860 12690 -790
rect 12760 -860 12800 -790
rect 12870 -860 12910 -790
rect 12980 -860 13020 -790
rect 13090 -860 13130 -790
rect 13200 -860 13240 -790
rect 13310 -860 13350 -790
rect 13420 -860 13460 -790
rect 13530 -860 13570 -790
rect 13640 -860 13680 -790
rect 13750 -860 13820 -790
rect 12220 -900 13820 -860
rect 12220 -970 12250 -900
rect 12320 -970 12360 -900
rect 12430 -970 12470 -900
rect 12540 -970 12580 -900
rect 12650 -970 12690 -900
rect 12760 -970 12800 -900
rect 12870 -970 12910 -900
rect 12980 -970 13020 -900
rect 13090 -970 13130 -900
rect 13200 -970 13240 -900
rect 13310 -970 13350 -900
rect 13420 -970 13460 -900
rect 13530 -970 13570 -900
rect 13640 -970 13680 -900
rect 13750 -970 13820 -900
rect 12220 -1020 13820 -970
rect 28700 -790 35790 -720
rect 35860 -790 35880 -720
rect 35950 -790 35970 -720
rect 36040 -790 36100 -720
rect 28700 -810 36100 -790
rect 28700 -880 35790 -810
rect 35860 -880 35880 -810
rect 35950 -880 35970 -810
rect 36040 -880 36100 -810
rect 28700 -900 36100 -880
rect 28700 -970 35790 -900
rect 35860 -970 35880 -900
rect 35950 -970 35970 -900
rect 36040 -970 36100 -900
rect 28700 -990 36100 -970
rect 28700 -1060 35790 -990
rect 35860 -1060 35880 -990
rect 35950 -1060 35970 -990
rect 36040 -1060 36100 -990
rect 28700 -1080 36100 -1060
rect 28700 -1150 35790 -1080
rect 35860 -1150 35880 -1080
rect 35950 -1150 35970 -1080
rect 36040 -1150 36100 -1080
rect 28700 -1170 36100 -1150
rect 28700 -1240 35790 -1170
rect 35860 -1240 35880 -1170
rect 35950 -1240 35970 -1170
rect 36040 -1240 36100 -1170
rect 28700 -1260 36100 -1240
rect 28700 -1330 35790 -1260
rect 35860 -1330 35880 -1260
rect 35950 -1330 35970 -1260
rect 36040 -1330 36100 -1260
rect 28700 -1350 36100 -1330
rect 28700 -1420 35790 -1350
rect 35860 -1420 35880 -1350
rect 35950 -1420 35970 -1350
rect 36040 -1420 36100 -1350
rect 28700 -1440 36100 -1420
rect 28700 -1510 35790 -1440
rect 35860 -1510 35880 -1440
rect 35950 -1510 35970 -1440
rect 36040 -1510 36100 -1440
rect 28700 -1530 36100 -1510
rect 28700 -1600 35790 -1530
rect 35860 -1600 35880 -1530
rect 35950 -1600 35970 -1530
rect 36040 -1600 36100 -1530
rect 28700 -1620 36100 -1600
rect 28700 -1690 35790 -1620
rect 35860 -1690 35880 -1620
rect 35950 -1690 35970 -1620
rect 36040 -1690 36100 -1620
rect 28700 -1710 36100 -1690
rect 28700 -1780 35790 -1710
rect 35860 -1780 35880 -1710
rect 35950 -1780 35970 -1710
rect 36040 -1780 36100 -1710
rect 28700 -1800 36100 -1780
rect 28700 -1870 35790 -1800
rect 35860 -1870 35880 -1800
rect 35950 -1870 35970 -1800
rect 36040 -1870 36100 -1800
rect 28700 -1890 36100 -1870
rect 28700 -1960 35790 -1890
rect 35860 -1960 35880 -1890
rect 35950 -1960 35970 -1890
rect 36040 -1960 36100 -1890
rect 28700 -1980 36100 -1960
rect 28700 -2050 35790 -1980
rect 35860 -2050 35880 -1980
rect 35950 -2050 35970 -1980
rect 36040 -2050 36100 -1980
rect 28700 -2070 36100 -2050
rect 28700 -2140 35790 -2070
rect 35860 -2140 35880 -2070
rect 35950 -2140 35970 -2070
rect 36040 -2140 36100 -2070
rect 28700 -2160 36100 -2140
rect 28700 -2230 35790 -2160
rect 35860 -2230 35880 -2160
rect 35950 -2230 35970 -2160
rect 36040 -2230 36100 -2160
rect 28700 -2250 36100 -2230
rect 28700 -2320 35790 -2250
rect 35860 -2320 35880 -2250
rect 35950 -2320 35970 -2250
rect 36040 -2320 36100 -2250
rect 28700 -2340 36100 -2320
rect 28700 -2410 35790 -2340
rect 35860 -2410 35880 -2340
rect 35950 -2410 35970 -2340
rect 36040 -2410 36100 -2340
rect 28700 -2430 36100 -2410
rect 28700 -2500 35790 -2430
rect 35860 -2500 35880 -2430
rect 35950 -2500 35970 -2430
rect 36040 -2500 36100 -2430
rect 28700 -2520 36100 -2500
rect 28700 -2590 35790 -2520
rect 35860 -2590 35880 -2520
rect 35950 -2590 35970 -2520
rect 36040 -2590 36100 -2520
rect 28700 -2610 36100 -2590
rect 28700 -2680 35790 -2610
rect 35860 -2680 35880 -2610
rect 35950 -2680 35970 -2610
rect 36040 -2680 36100 -2610
rect 28700 -2700 36100 -2680
rect 11760 -2780 13360 -2730
rect 11760 -2850 11790 -2780
rect 11860 -2850 11900 -2780
rect 11970 -2850 12010 -2780
rect 12080 -2850 12120 -2780
rect 12190 -2850 12230 -2780
rect 12300 -2850 12340 -2780
rect 12410 -2850 12450 -2780
rect 12520 -2850 12560 -2780
rect 12630 -2850 12670 -2780
rect 12740 -2850 12780 -2780
rect 12850 -2850 12890 -2780
rect 12960 -2850 13000 -2780
rect 13070 -2850 13110 -2780
rect 13180 -2850 13220 -2780
rect 13290 -2850 13360 -2780
rect 11760 -2890 13360 -2850
rect 11760 -2960 11790 -2890
rect 11860 -2960 11900 -2890
rect 11970 -2960 12010 -2890
rect 12080 -2960 12120 -2890
rect 12190 -2960 12230 -2890
rect 12300 -2960 12340 -2890
rect 12410 -2960 12450 -2890
rect 12520 -2960 12560 -2890
rect 12630 -2960 12670 -2890
rect 12740 -2960 12780 -2890
rect 12850 -2960 12890 -2890
rect 12960 -2960 13000 -2890
rect 13070 -2960 13110 -2890
rect 13180 -2960 13220 -2890
rect 13290 -2960 13360 -2890
rect 11760 -2990 13360 -2960
rect 28700 -2770 35790 -2700
rect 35860 -2770 35880 -2700
rect 35950 -2770 35970 -2700
rect 36040 -2770 36100 -2700
rect 28700 -2790 36100 -2770
rect 28700 -2860 35790 -2790
rect 35860 -2860 35880 -2790
rect 35950 -2860 35970 -2790
rect 36040 -2860 36100 -2790
rect 28700 -2880 36100 -2860
rect 28700 -2950 35790 -2880
rect 35860 -2950 35880 -2880
rect 35950 -2950 35970 -2880
rect 36040 -2950 36100 -2880
rect 28700 -2970 36100 -2950
rect 22320 -3050 22650 -3030
rect 22320 -3120 22340 -3050
rect 22410 -3120 22450 -3050
rect 22520 -3120 22560 -3050
rect 22630 -3120 22650 -3050
rect 22320 -3160 22650 -3120
rect 22320 -3230 22340 -3160
rect 22410 -3230 22450 -3160
rect 22520 -3230 22560 -3160
rect 22630 -3230 22650 -3160
rect 22320 -3270 22650 -3230
rect 22320 -3340 22340 -3270
rect 22410 -3340 22450 -3270
rect 22520 -3340 22560 -3270
rect 22630 -3340 22650 -3270
rect 22320 -3360 22650 -3340
rect 28700 -3040 35790 -2970
rect 35860 -3040 35880 -2970
rect 35950 -3040 35970 -2970
rect 36040 -3040 36100 -2970
rect 28700 -3060 36100 -3040
rect 28700 -3130 35790 -3060
rect 35860 -3130 35880 -3060
rect 35950 -3130 35970 -3060
rect 36040 -3130 36100 -3060
rect 28700 -3150 36100 -3130
rect 28700 -3220 35790 -3150
rect 35860 -3220 35880 -3150
rect 35950 -3220 35970 -3150
rect 36040 -3220 36100 -3150
rect 28700 -3240 36100 -3220
rect 28700 -3310 35790 -3240
rect 35860 -3310 35880 -3240
rect 35950 -3310 35970 -3240
rect 36040 -3310 36100 -3240
rect 28700 -3330 36100 -3310
rect 28700 -3400 35790 -3330
rect 35860 -3400 35880 -3330
rect 35950 -3400 35970 -3330
rect 36040 -3400 36100 -3330
rect 28700 -3460 36100 -3400
rect 28700 -3530 35790 -3460
rect 35860 -3530 35880 -3460
rect 35950 -3530 35970 -3460
rect 36040 -3530 36100 -3460
rect 28700 -3550 36100 -3530
rect 28700 -3620 35790 -3550
rect 35860 -3620 35880 -3550
rect 35950 -3620 35970 -3550
rect 36040 -3620 36100 -3550
rect 28700 -3640 36100 -3620
rect 20020 -3690 20500 -3660
rect 20020 -3760 20070 -3690
rect 20140 -3760 20180 -3690
rect 20250 -3760 20290 -3690
rect 20360 -3760 20400 -3690
rect 20470 -3760 20500 -3690
rect 20020 -3800 20500 -3760
rect 20020 -3870 20070 -3800
rect 20140 -3870 20180 -3800
rect 20250 -3870 20290 -3800
rect 20360 -3870 20400 -3800
rect 20470 -3870 20500 -3800
rect 20020 -3920 20500 -3870
rect 24500 -3690 24980 -3660
rect 24500 -3760 24550 -3690
rect 24620 -3760 24660 -3690
rect 24730 -3760 24770 -3690
rect 24840 -3760 24880 -3690
rect 24950 -3760 24980 -3690
rect 24500 -3800 24980 -3760
rect 24500 -3870 24550 -3800
rect 24620 -3870 24660 -3800
rect 24730 -3870 24770 -3800
rect 24840 -3870 24880 -3800
rect 24950 -3870 24980 -3800
rect 24500 -3920 24980 -3870
rect 28700 -3710 35790 -3640
rect 35860 -3710 35880 -3640
rect 35950 -3710 35970 -3640
rect 36040 -3710 36100 -3640
rect 28700 -3730 36100 -3710
rect 28700 -3800 35790 -3730
rect 35860 -3800 35880 -3730
rect 35950 -3800 35970 -3730
rect 36040 -3800 36100 -3730
rect 28700 -3820 36100 -3800
rect 28700 -3890 35790 -3820
rect 35860 -3890 35880 -3820
rect 35950 -3890 35970 -3820
rect 36040 -3890 36100 -3820
rect 28700 -3910 36100 -3890
rect 8180 -6220 8200 -6150
rect 8270 -6220 8300 -6150
rect 8370 -6220 8400 -6150
rect 8470 -6220 8490 -6150
rect 8180 -6250 8490 -6220
rect 8180 -6320 8200 -6250
rect 8270 -6320 8300 -6250
rect 8370 -6320 8400 -6250
rect 8470 -6320 8490 -6250
rect 8180 -6420 8490 -6320
rect 6440 -6460 7340 -6420
rect 6440 -6520 7050 -6460
rect 7110 -6520 7150 -6460
rect 7210 -6520 7250 -6460
rect 7310 -6520 7340 -6460
rect 6440 -6560 7340 -6520
rect 6440 -6620 7050 -6560
rect 7110 -6620 7150 -6560
rect 7210 -6620 7250 -6560
rect 7310 -6620 7340 -6560
rect -640 -6670 6190 -6640
rect -640 -6680 4770 -6670
rect -880 -6720 4770 -6680
rect -880 -6790 -840 -6720
rect -770 -6790 -710 -6720
rect -640 -6730 4770 -6720
rect 4830 -6730 4870 -6670
rect 4930 -6730 4970 -6670
rect 5030 -6730 6190 -6670
rect -640 -6770 6190 -6730
rect -640 -6790 4770 -6770
rect -880 -6830 4770 -6790
rect 4830 -6830 4870 -6770
rect 4930 -6830 4970 -6770
rect 5030 -6830 6190 -6770
rect -880 -6900 -840 -6830
rect -770 -6900 -710 -6830
rect -640 -6870 6190 -6830
rect 6440 -6660 7340 -6620
rect 6440 -6720 7050 -6660
rect 7110 -6720 7150 -6660
rect 7210 -6720 7250 -6660
rect 7310 -6720 7340 -6660
rect 6440 -6760 7340 -6720
rect 6440 -6820 7050 -6760
rect 7110 -6820 7150 -6760
rect 7210 -6820 7250 -6760
rect 7310 -6820 7340 -6760
rect 6440 -6850 7340 -6820
rect 7560 -6460 8490 -6420
rect 28700 -3980 35790 -3910
rect 35860 -3980 35880 -3910
rect 35950 -3980 35970 -3910
rect 36040 -3980 36100 -3910
rect 28700 -4000 36100 -3980
rect 28700 -4070 35790 -4000
rect 35860 -4070 35880 -4000
rect 35950 -4070 35970 -4000
rect 36040 -4070 36100 -4000
rect 28700 -4090 36100 -4070
rect 28700 -4160 35790 -4090
rect 35860 -4160 35880 -4090
rect 35950 -4160 35970 -4090
rect 36040 -4160 36100 -4090
rect 28700 -4180 36100 -4160
rect 28700 -4250 35790 -4180
rect 35860 -4250 35880 -4180
rect 35950 -4250 35970 -4180
rect 36040 -4250 36100 -4180
rect 28700 -4270 36100 -4250
rect 28700 -4340 35790 -4270
rect 35860 -4340 35880 -4270
rect 35950 -4340 35970 -4270
rect 36040 -4340 36100 -4270
rect 28700 -4360 36100 -4340
rect 28700 -4430 35790 -4360
rect 35860 -4430 35880 -4360
rect 35950 -4430 35970 -4360
rect 36040 -4430 36100 -4360
rect 28700 -4450 36100 -4430
rect 28700 -4520 35790 -4450
rect 35860 -4520 35880 -4450
rect 35950 -4520 35970 -4450
rect 36040 -4520 36100 -4450
rect 28700 -4540 36100 -4520
rect 28700 -4610 35790 -4540
rect 35860 -4610 35880 -4540
rect 35950 -4610 35970 -4540
rect 36040 -4610 36100 -4540
rect 28700 -4630 36100 -4610
rect 28700 -4700 35790 -4630
rect 35860 -4700 35880 -4630
rect 35950 -4700 35970 -4630
rect 36040 -4700 36100 -4630
rect 28700 -4720 36100 -4700
rect 28700 -4790 35790 -4720
rect 35860 -4790 35880 -4720
rect 35950 -4790 35970 -4720
rect 36040 -4790 36100 -4720
rect 28700 -4810 36100 -4790
rect 28700 -4880 35790 -4810
rect 35860 -4880 35880 -4810
rect 35950 -4880 35970 -4810
rect 36040 -4880 36100 -4810
rect 28700 -4900 36100 -4880
rect 28700 -4970 35790 -4900
rect 35860 -4970 35880 -4900
rect 35950 -4970 35970 -4900
rect 36040 -4970 36100 -4900
rect 28700 -4990 36100 -4970
rect 28700 -5060 35790 -4990
rect 35860 -5060 35880 -4990
rect 35950 -5060 35970 -4990
rect 36040 -5060 36100 -4990
rect 28700 -5080 36100 -5060
rect 28700 -5150 35790 -5080
rect 35860 -5150 35880 -5080
rect 35950 -5150 35970 -5080
rect 36040 -5150 36100 -5080
rect 28700 -5170 36100 -5150
rect 28700 -5240 35790 -5170
rect 35860 -5240 35880 -5170
rect 35950 -5240 35970 -5170
rect 36040 -5240 36100 -5170
rect 28700 -5260 36100 -5240
rect 28700 -5330 35790 -5260
rect 35860 -5330 35880 -5260
rect 35950 -5330 35970 -5260
rect 36040 -5330 36100 -5260
rect 28700 -5350 36100 -5330
rect 28700 -5420 35790 -5350
rect 35860 -5420 35880 -5350
rect 35950 -5420 35970 -5350
rect 36040 -5420 36100 -5350
rect 28700 -5440 36100 -5420
rect 28700 -5510 35790 -5440
rect 35860 -5510 35880 -5440
rect 35950 -5510 35970 -5440
rect 36040 -5510 36100 -5440
rect 28700 -5530 36100 -5510
rect 28700 -5600 35790 -5530
rect 35860 -5600 35880 -5530
rect 35950 -5600 35970 -5530
rect 36040 -5600 36100 -5530
rect 28700 -5620 36100 -5600
rect 28700 -5690 35790 -5620
rect 35860 -5690 35880 -5620
rect 35950 -5690 35970 -5620
rect 36040 -5690 36100 -5620
rect 28700 -5710 36100 -5690
rect 28700 -5780 35790 -5710
rect 35860 -5780 35880 -5710
rect 35950 -5780 35970 -5710
rect 36040 -5780 36100 -5710
rect 28700 -5800 36100 -5780
rect 28700 -5870 35790 -5800
rect 35860 -5870 35880 -5800
rect 35950 -5870 35970 -5800
rect 36040 -5870 36100 -5800
rect 28700 -5890 36100 -5870
rect 28700 -5960 35790 -5890
rect 35860 -5960 35880 -5890
rect 35950 -5960 35970 -5890
rect 36040 -5960 36100 -5890
rect 28700 -5980 36100 -5960
rect 28700 -6050 35790 -5980
rect 35860 -6050 35880 -5980
rect 35950 -6050 35970 -5980
rect 36040 -6050 36100 -5980
rect 28700 -6070 36100 -6050
rect 28700 -6140 35790 -6070
rect 35860 -6140 35880 -6070
rect 35950 -6140 35970 -6070
rect 36040 -6140 36100 -6070
rect 28700 -6160 36100 -6140
rect 28700 -6230 35790 -6160
rect 35860 -6230 35880 -6160
rect 35950 -6230 35970 -6160
rect 36040 -6230 36100 -6160
rect 28700 -6250 36100 -6230
rect 28700 -6320 35790 -6250
rect 35860 -6320 35880 -6250
rect 35950 -6320 35970 -6250
rect 36040 -6320 36100 -6250
rect 28700 -6340 36100 -6320
rect 28700 -6410 35790 -6340
rect 35860 -6410 35880 -6340
rect 35950 -6410 35970 -6340
rect 36040 -6410 36100 -6340
rect 28700 -6450 36100 -6410
rect 7560 -6520 7590 -6460
rect 7650 -6520 7690 -6460
rect 7750 -6520 7790 -6460
rect 7850 -6520 8490 -6460
rect 7560 -6560 8490 -6520
rect 7560 -6620 7590 -6560
rect 7650 -6620 7690 -6560
rect 7750 -6620 7790 -6560
rect 7850 -6620 8490 -6560
rect 7560 -6660 8490 -6620
rect 15380 -6500 15660 -6470
rect 15380 -6570 15420 -6500
rect 15490 -6570 15550 -6500
rect 15620 -6570 15660 -6500
rect 15380 -6610 15660 -6570
rect 15380 -6640 15420 -6610
rect 7560 -6720 7590 -6660
rect 7650 -6720 7690 -6660
rect 7750 -6720 7790 -6660
rect 7850 -6720 8490 -6660
rect 7560 -6760 8490 -6720
rect 7560 -6820 7590 -6760
rect 7650 -6820 7690 -6760
rect 7750 -6820 7790 -6760
rect 7850 -6820 8490 -6760
rect 7560 -6850 8490 -6820
rect 8710 -6670 15420 -6640
rect 8710 -6730 9870 -6670
rect 9930 -6730 9970 -6670
rect 10030 -6730 10070 -6670
rect 10130 -6680 15420 -6670
rect 15490 -6680 15550 -6610
rect 15620 -6680 15660 -6610
rect 10130 -6720 15660 -6680
rect 10130 -6730 15420 -6720
rect 8710 -6770 15420 -6730
rect 8710 -6830 9870 -6770
rect 9930 -6830 9970 -6770
rect 10030 -6830 10070 -6770
rect 10130 -6790 15420 -6770
rect 15490 -6790 15550 -6720
rect 15620 -6790 15660 -6720
rect 10130 -6830 15660 -6790
rect -640 -6900 4770 -6870
rect -880 -6930 4770 -6900
rect 4830 -6930 4870 -6870
rect 4930 -6930 4970 -6870
rect 5030 -6930 6190 -6870
rect -880 -6950 6190 -6930
rect -1860 -7630 150 -7450
rect -1860 -7700 -160 -7630
rect -90 -7700 -70 -7630
rect 0 -7700 20 -7630
rect 90 -7700 150 -7630
rect -1860 -7720 150 -7700
rect -1860 -7790 -160 -7720
rect -90 -7790 -70 -7720
rect 0 -7790 20 -7720
rect 90 -7790 150 -7720
rect -1860 -7810 150 -7790
rect -2220 -7870 -2000 -7850
rect -2220 -7940 -2200 -7870
rect -2130 -7940 -2090 -7870
rect -2020 -7940 -2000 -7870
rect -2220 -7980 -2000 -7940
rect -2220 -8050 -2200 -7980
rect -2130 -8050 -2090 -7980
rect -2020 -8050 -2000 -7980
rect -2220 -8090 -2000 -8050
rect -2220 -8160 -2200 -8090
rect -2130 -8160 -2090 -8090
rect -2020 -8160 -2000 -8090
rect -2220 -8200 -2000 -8160
rect -2220 -8270 -2200 -8200
rect -2130 -8270 -2090 -8200
rect -2020 -8270 -2000 -8200
rect -2220 -8290 -2000 -8270
rect -1860 -7880 -160 -7810
rect -90 -7880 -70 -7810
rect 0 -7880 20 -7810
rect 90 -7880 150 -7810
rect -1860 -7900 150 -7880
rect -1860 -7970 -160 -7900
rect -90 -7970 -70 -7900
rect 0 -7970 20 -7900
rect 90 -7970 150 -7900
rect -1860 -7990 150 -7970
rect -1860 -8060 -160 -7990
rect -90 -8060 -70 -7990
rect 0 -8060 20 -7990
rect 90 -8060 150 -7990
rect -1860 -8080 150 -8060
rect -1860 -8150 -160 -8080
rect -90 -8150 -70 -8080
rect 0 -8150 20 -8080
rect 90 -8150 150 -8080
rect -1860 -8170 150 -8150
rect -1860 -8240 -160 -8170
rect -90 -8240 -70 -8170
rect 0 -8240 20 -8170
rect 90 -8240 150 -8170
rect -1860 -8260 150 -8240
rect -1860 -8330 -160 -8260
rect -90 -8330 -70 -8260
rect 0 -8330 20 -8260
rect 90 -8330 150 -8260
rect -1860 -8350 150 -8330
rect -1860 -8420 -160 -8350
rect -90 -8420 -70 -8350
rect 0 -8420 20 -8350
rect 90 -8420 150 -8350
rect -1860 -8440 150 -8420
rect -1860 -8510 -160 -8440
rect -90 -8510 -70 -8440
rect 0 -8510 20 -8440
rect 90 -8510 150 -8440
rect -1860 -8530 150 -8510
rect -1860 -8600 -160 -8530
rect -90 -8600 -70 -8530
rect 0 -8600 20 -8530
rect 90 -8600 150 -8530
rect -1860 -8620 150 -8600
rect -2160 -8640 -1940 -8620
rect -2160 -8710 -2140 -8640
rect -2070 -8710 -2030 -8640
rect -1960 -8710 -1940 -8640
rect -2160 -8750 -1940 -8710
rect -2160 -8820 -2140 -8750
rect -2070 -8820 -2030 -8750
rect -1960 -8820 -1940 -8750
rect -2160 -8860 -1940 -8820
rect -2160 -8930 -2140 -8860
rect -2070 -8930 -2030 -8860
rect -1960 -8930 -1940 -8860
rect -2160 -8970 -1940 -8930
rect -2160 -9040 -2140 -8970
rect -2070 -9040 -2030 -8970
rect -1960 -9040 -1940 -8970
rect -2160 -9060 -1940 -9040
rect -1860 -8690 -160 -8620
rect -90 -8690 -70 -8620
rect 0 -8690 20 -8620
rect 90 -8690 150 -8620
rect -1860 -8710 150 -8690
rect -1860 -8780 -160 -8710
rect -90 -8780 -70 -8710
rect 0 -8780 20 -8710
rect 90 -8780 150 -8710
rect -1860 -8800 150 -8780
rect -1860 -8870 -160 -8800
rect -90 -8870 -70 -8800
rect 0 -8870 20 -8800
rect 90 -8870 150 -8800
rect -1860 -9060 150 -8870
rect 5880 -9620 6190 -6950
rect -270 -9660 6190 -9620
rect -270 -9730 -240 -9660
rect -170 -9730 -130 -9660
rect -60 -9730 -20 -9660
rect 50 -9730 90 -9660
rect 160 -9730 6190 -9660
rect -270 -9790 6190 -9730
rect -270 -9860 -240 -9790
rect -170 -9860 -130 -9790
rect -60 -9860 -20 -9790
rect 50 -9860 90 -9790
rect 160 -9860 6190 -9790
rect -270 -9900 6190 -9860
rect 1080 -10340 2680 -10310
rect 1080 -10410 1150 -10340
rect 1220 -10410 1260 -10340
rect 1330 -10410 1370 -10340
rect 1440 -10410 1480 -10340
rect 1550 -10410 1590 -10340
rect 1660 -10410 1700 -10340
rect 1770 -10410 1810 -10340
rect 1880 -10410 1920 -10340
rect 1990 -10410 2030 -10340
rect 2100 -10410 2140 -10340
rect 2210 -10410 2250 -10340
rect 2320 -10410 2360 -10340
rect 2430 -10410 2470 -10340
rect 2540 -10410 2580 -10340
rect 2650 -10410 2680 -10340
rect 1080 -10450 2680 -10410
rect 1080 -10520 1150 -10450
rect 1220 -10520 1260 -10450
rect 1330 -10520 1370 -10450
rect 1440 -10520 1480 -10450
rect 1550 -10520 1590 -10450
rect 1660 -10520 1700 -10450
rect 1770 -10520 1810 -10450
rect 1880 -10520 1920 -10450
rect 1990 -10520 2030 -10450
rect 2100 -10520 2140 -10450
rect 2210 -10520 2250 -10450
rect 2320 -10520 2360 -10450
rect 2430 -10520 2470 -10450
rect 2540 -10520 2580 -10450
rect 2650 -10520 2680 -10450
rect 1080 -10570 2680 -10520
rect 2210 -12300 3810 -12250
rect 2210 -12370 2240 -12300
rect 2310 -12370 2350 -12300
rect 2420 -12370 2460 -12300
rect 2530 -12370 2570 -12300
rect 2640 -12370 2680 -12300
rect 2750 -12370 2790 -12300
rect 2860 -12370 2900 -12300
rect 2970 -12370 3010 -12300
rect 3080 -12370 3120 -12300
rect 3190 -12370 3230 -12300
rect 3300 -12370 3340 -12300
rect 3410 -12370 3450 -12300
rect 3520 -12370 3560 -12300
rect 3630 -12370 3670 -12300
rect 3740 -12370 3810 -12300
rect 2210 -12410 3810 -12370
rect 2210 -12480 2240 -12410
rect 2310 -12480 2350 -12410
rect 2420 -12480 2460 -12410
rect 2530 -12480 2570 -12410
rect 2640 -12480 2680 -12410
rect 2750 -12480 2790 -12410
rect 2860 -12480 2900 -12410
rect 2970 -12480 3010 -12410
rect 3080 -12480 3120 -12410
rect 3190 -12480 3230 -12410
rect 3300 -12480 3340 -12410
rect 3410 -12480 3450 -12410
rect 3520 -12480 3560 -12410
rect 3630 -12480 3670 -12410
rect 3740 -12480 3810 -12410
rect 2210 -12510 3810 -12480
rect 5880 -13220 6190 -9900
rect 8710 -6870 15420 -6830
rect 8710 -6930 9870 -6870
rect 9930 -6930 9970 -6870
rect 10030 -6930 10070 -6870
rect 10130 -6900 15420 -6870
rect 15490 -6900 15550 -6830
rect 15620 -6900 15660 -6830
rect 10130 -6930 15660 -6900
rect 8710 -6950 15660 -6930
rect 8710 -8250 9020 -6950
rect 8710 -8320 8730 -8250
rect 8800 -8320 8830 -8250
rect 8900 -8320 8930 -8250
rect 9000 -8320 9020 -8250
rect 8710 -8350 9020 -8320
rect 8710 -8420 8730 -8350
rect 8800 -8420 8830 -8350
rect 8900 -8420 8930 -8350
rect 9000 -8420 9020 -8350
rect 8710 -9620 9020 -8420
rect 14590 -8230 14900 -8210
rect 14590 -8300 14600 -8230
rect 14670 -8300 14700 -8230
rect 14770 -8300 14810 -8230
rect 14880 -8300 14900 -8230
rect 14590 -8340 14900 -8300
rect 14590 -8410 14600 -8340
rect 14670 -8410 14700 -8340
rect 14770 -8410 14810 -8340
rect 14880 -8410 14900 -8340
rect 14590 -8450 14900 -8410
rect 14590 -8520 14600 -8450
rect 14670 -8520 14700 -8450
rect 14770 -8520 14810 -8450
rect 14880 -8520 14900 -8450
rect 14590 -8540 14900 -8520
rect 19210 -8560 19530 -8530
rect 19210 -8630 19230 -8560
rect 19300 -8630 19330 -8560
rect 19400 -8630 19430 -8560
rect 19500 -8630 19530 -8560
rect 19210 -8660 19530 -8630
rect 19210 -8730 19230 -8660
rect 19300 -8730 19330 -8660
rect 19400 -8730 19430 -8660
rect 19500 -8730 19530 -8660
rect 19210 -8760 19530 -8730
rect 19210 -8830 19230 -8760
rect 19300 -8830 19330 -8760
rect 19400 -8830 19430 -8760
rect 19500 -8830 19530 -8760
rect 19210 -8850 19530 -8830
rect 19940 -9000 20260 -8970
rect 19940 -9070 19960 -9000
rect 20030 -9070 20060 -9000
rect 20130 -9070 20160 -9000
rect 20230 -9070 20260 -9000
rect 19940 -9100 20260 -9070
rect 19940 -9170 19960 -9100
rect 20030 -9170 20060 -9100
rect 20130 -9170 20160 -9100
rect 20230 -9170 20260 -9100
rect 19940 -9200 20260 -9170
rect 19940 -9270 19960 -9200
rect 20030 -9270 20060 -9200
rect 20130 -9270 20160 -9200
rect 20230 -9270 20260 -9200
rect 19940 -9290 20260 -9270
rect 8710 -9660 15170 -9620
rect 8710 -9730 14720 -9660
rect 14790 -9730 14830 -9660
rect 14900 -9730 14940 -9660
rect 15010 -9730 15050 -9660
rect 15120 -9730 15170 -9660
rect 8710 -9790 15170 -9730
rect 8710 -9860 14720 -9790
rect 14790 -9860 14830 -9790
rect 14900 -9860 14940 -9790
rect 15010 -9860 15050 -9790
rect 15120 -9860 15170 -9790
rect 8710 -9900 15170 -9860
rect 8710 -13220 9020 -9900
rect 12220 -10370 13820 -10340
rect 12220 -10440 12290 -10370
rect 12360 -10440 12400 -10370
rect 12470 -10440 12510 -10370
rect 12580 -10440 12620 -10370
rect 12690 -10440 12730 -10370
rect 12800 -10440 12840 -10370
rect 12910 -10440 12950 -10370
rect 13020 -10440 13060 -10370
rect 13130 -10440 13170 -10370
rect 13240 -10440 13280 -10370
rect 13350 -10440 13390 -10370
rect 13460 -10440 13500 -10370
rect 13570 -10440 13610 -10370
rect 13680 -10440 13720 -10370
rect 13790 -10440 13820 -10370
rect 12220 -10480 13820 -10440
rect 12220 -10550 12290 -10480
rect 12360 -10550 12400 -10480
rect 12470 -10550 12510 -10480
rect 12580 -10550 12620 -10480
rect 12690 -10550 12730 -10480
rect 12800 -10550 12840 -10480
rect 12910 -10550 12950 -10480
rect 13020 -10550 13060 -10480
rect 13130 -10550 13170 -10480
rect 13240 -10550 13280 -10480
rect 13350 -10550 13390 -10480
rect 13460 -10550 13500 -10480
rect 13570 -10550 13610 -10480
rect 13680 -10550 13720 -10480
rect 13790 -10550 13820 -10480
rect 12220 -10600 13820 -10550
rect 11090 -12300 12690 -12250
rect 11090 -12370 11120 -12300
rect 11190 -12370 11230 -12300
rect 11300 -12370 11340 -12300
rect 11410 -12370 11450 -12300
rect 11520 -12370 11560 -12300
rect 11630 -12370 11670 -12300
rect 11740 -12370 11780 -12300
rect 11850 -12370 11890 -12300
rect 11960 -12370 12000 -12300
rect 12070 -12370 12110 -12300
rect 12180 -12370 12220 -12300
rect 12290 -12370 12330 -12300
rect 12400 -12370 12440 -12300
rect 12510 -12370 12550 -12300
rect 12620 -12370 12690 -12300
rect 11090 -12410 12690 -12370
rect 11090 -12480 11120 -12410
rect 11190 -12480 11230 -12410
rect 11300 -12480 11340 -12410
rect 11410 -12480 11450 -12410
rect 11520 -12480 11560 -12410
rect 11630 -12480 11670 -12410
rect 11740 -12480 11780 -12410
rect 11850 -12480 11890 -12410
rect 11960 -12480 12000 -12410
rect 12070 -12480 12110 -12410
rect 12180 -12480 12220 -12410
rect 12290 -12480 12330 -12410
rect 12400 -12480 12440 -12410
rect 12510 -12480 12550 -12410
rect 12620 -12480 12690 -12410
rect 11090 -12510 12690 -12480
rect 5880 -13250 7310 -13220
rect 5880 -13310 7010 -13250
rect 7070 -13310 7110 -13250
rect 7170 -13310 7210 -13250
rect 7270 -13310 7310 -13250
rect 5880 -13340 7310 -13310
rect 5880 -13400 7010 -13340
rect 7070 -13400 7110 -13340
rect 7170 -13400 7210 -13340
rect 7270 -13400 7310 -13340
rect 5880 -13430 7310 -13400
rect 5880 -13490 7010 -13430
rect 7070 -13490 7110 -13430
rect 7170 -13490 7210 -13430
rect 7270 -13490 7310 -13430
rect 5880 -13530 7310 -13490
rect 5880 -13590 7010 -13530
rect 7070 -13590 7110 -13530
rect 7170 -13590 7210 -13530
rect 7270 -13590 7310 -13530
rect 5880 -13620 7310 -13590
rect 5880 -13680 7010 -13620
rect 7070 -13680 7110 -13620
rect 7170 -13680 7210 -13620
rect 7270 -13680 7310 -13620
rect 5880 -13710 7310 -13680
rect 5880 -13770 7010 -13710
rect 7070 -13770 7110 -13710
rect 7170 -13770 7210 -13710
rect 7270 -13770 7310 -13710
rect 5880 -13800 7310 -13770
rect 7590 -13250 9020 -13220
rect 7590 -13310 7630 -13250
rect 7690 -13310 7730 -13250
rect 7790 -13310 7830 -13250
rect 7890 -13310 9020 -13250
rect 7590 -13340 9020 -13310
rect 7590 -13400 7630 -13340
rect 7690 -13400 7730 -13340
rect 7790 -13400 7830 -13340
rect 7890 -13400 9020 -13340
rect 7590 -13430 9020 -13400
rect 7590 -13490 7630 -13430
rect 7690 -13490 7730 -13430
rect 7790 -13490 7830 -13430
rect 7890 -13490 9020 -13430
rect 7590 -13530 9020 -13490
rect 7590 -13590 7630 -13530
rect 7690 -13590 7730 -13530
rect 7790 -13590 7830 -13530
rect 7890 -13590 9020 -13530
rect 7590 -13620 9020 -13590
rect 7590 -13680 7630 -13620
rect 7690 -13680 7730 -13620
rect 7790 -13680 7830 -13620
rect 7890 -13680 9020 -13620
rect 7590 -13710 9020 -13680
rect 7590 -13770 7630 -13710
rect 7690 -13770 7730 -13710
rect 7790 -13770 7830 -13710
rect 7890 -13770 9020 -13710
rect 7590 -13800 9020 -13770
rect 19210 -14220 19530 -14190
rect 19210 -14290 19230 -14220
rect 19300 -14290 19330 -14220
rect 19400 -14290 19430 -14220
rect 19500 -14290 19530 -14220
rect 19210 -14320 19530 -14290
rect 19210 -14390 19230 -14320
rect 19300 -14390 19330 -14320
rect 19400 -14390 19430 -14320
rect 19500 -14390 19530 -14320
rect 19210 -14420 19530 -14390
rect 19210 -14490 19230 -14420
rect 19300 -14490 19330 -14420
rect 19400 -14490 19430 -14420
rect 19500 -14490 19530 -14420
rect 19210 -14510 19530 -14490
rect 20460 -14870 20780 -14840
rect 20460 -14940 20480 -14870
rect 20550 -14940 20580 -14870
rect 20650 -14940 20680 -14870
rect 20750 -14940 20780 -14870
rect 20460 -14970 20780 -14940
rect 20460 -15040 20480 -14970
rect 20550 -15040 20580 -14970
rect 20650 -15040 20680 -14970
rect 20750 -15040 20780 -14970
rect 20460 -15070 20780 -15040
rect 20460 -15140 20480 -15070
rect 20550 -15140 20580 -15070
rect 20650 -15140 20680 -15070
rect 20750 -15140 20780 -15070
rect 20460 -15160 20780 -15140
rect 5010 -17100 5330 -17070
rect 5010 -17160 5040 -17100
rect 5100 -17160 5140 -17100
rect 5200 -17160 5240 -17100
rect 5300 -17160 5330 -17100
rect 5010 -17200 5330 -17160
rect 5010 -17260 5040 -17200
rect 5100 -17260 5140 -17200
rect 5200 -17260 5240 -17200
rect 5300 -17260 5330 -17200
rect 5010 -17300 5330 -17260
rect 5010 -17360 5040 -17300
rect 5100 -17360 5140 -17300
rect 5200 -17360 5240 -17300
rect 5300 -17360 5330 -17300
rect 2210 -22660 3810 -22630
rect 2210 -22730 2280 -22660
rect 2350 -22730 2390 -22660
rect 2460 -22730 2500 -22660
rect 2570 -22730 2610 -22660
rect 2680 -22730 2720 -22660
rect 2790 -22730 2830 -22660
rect 2900 -22730 2940 -22660
rect 3010 -22730 3050 -22660
rect 3120 -22730 3160 -22660
rect 3230 -22730 3270 -22660
rect 3340 -22730 3380 -22660
rect 3450 -22730 3490 -22660
rect 3560 -22730 3600 -22660
rect 3670 -22730 3710 -22660
rect 3780 -22730 3810 -22660
rect 2210 -22770 3810 -22730
rect 2210 -22840 2280 -22770
rect 2350 -22840 2390 -22770
rect 2460 -22840 2500 -22770
rect 2570 -22840 2610 -22770
rect 2680 -22840 2720 -22770
rect 2790 -22840 2830 -22770
rect 2900 -22840 2940 -22770
rect 3010 -22840 3050 -22770
rect 3120 -22840 3160 -22770
rect 3230 -22840 3270 -22770
rect 3340 -22840 3380 -22770
rect 3450 -22840 3490 -22770
rect 3560 -22840 3600 -22770
rect 3670 -22840 3710 -22770
rect 3780 -22840 3810 -22770
rect 2210 -22890 3810 -22840
rect 5010 -23690 5330 -17360
rect 9570 -17100 9890 -17070
rect 9570 -17160 9600 -17100
rect 9660 -17160 9700 -17100
rect 9760 -17160 9800 -17100
rect 9860 -17160 9890 -17100
rect 9570 -17200 9890 -17160
rect 9570 -17260 9600 -17200
rect 9660 -17260 9700 -17200
rect 9760 -17260 9800 -17200
rect 9860 -17260 9890 -17200
rect 9570 -17300 9890 -17260
rect 9570 -17360 9600 -17300
rect 9660 -17360 9700 -17300
rect 9760 -17360 9800 -17300
rect 9860 -17360 9890 -17300
rect 7210 -17600 7650 -17580
rect 7210 -17670 7230 -17600
rect 7300 -17670 7340 -17600
rect 7410 -17670 7450 -17600
rect 7520 -17670 7560 -17600
rect 7630 -17670 7650 -17600
rect 7210 -17710 7650 -17670
rect 7210 -17780 7230 -17710
rect 7300 -17780 7340 -17710
rect 7410 -17780 7450 -17710
rect 7520 -17780 7560 -17710
rect 7630 -17780 7650 -17710
rect 7210 -17820 7650 -17780
rect 7210 -17890 7230 -17820
rect 7300 -17890 7340 -17820
rect 7410 -17890 7450 -17820
rect 7520 -17890 7560 -17820
rect 7630 -17890 7650 -17820
rect 7210 -17930 7650 -17890
rect 7210 -18000 7230 -17930
rect 7300 -18000 7340 -17930
rect 7410 -18000 7450 -17930
rect 7520 -18000 7560 -17930
rect 7630 -18000 7650 -17930
rect 7210 -18020 7650 -18000
rect 9570 -23690 9890 -17360
rect 19210 -20290 19530 -20260
rect 19210 -20360 19230 -20290
rect 19300 -20360 19330 -20290
rect 19400 -20360 19430 -20290
rect 19500 -20360 19530 -20290
rect 19210 -20390 19530 -20360
rect 19210 -20460 19230 -20390
rect 19300 -20460 19330 -20390
rect 19400 -20460 19430 -20390
rect 19500 -20460 19530 -20390
rect 19210 -20490 19530 -20460
rect 19210 -20560 19230 -20490
rect 19300 -20560 19330 -20490
rect 19400 -20560 19430 -20490
rect 19500 -20560 19530 -20490
rect 19210 -20580 19530 -20560
rect 20020 -20720 20340 -20690
rect 20020 -20790 20040 -20720
rect 20110 -20790 20140 -20720
rect 20210 -20790 20240 -20720
rect 20310 -20790 20340 -20720
rect 20020 -20820 20340 -20790
rect 20020 -20890 20040 -20820
rect 20110 -20890 20140 -20820
rect 20210 -20890 20240 -20820
rect 20310 -20890 20340 -20820
rect 20020 -20920 20340 -20890
rect 20020 -20990 20040 -20920
rect 20110 -20990 20140 -20920
rect 20210 -20990 20240 -20920
rect 20310 -20990 20340 -20920
rect 20020 -21010 20340 -20990
rect 11090 -22660 12690 -22630
rect 11090 -22730 11160 -22660
rect 11230 -22730 11270 -22660
rect 11340 -22730 11380 -22660
rect 11450 -22730 11490 -22660
rect 11560 -22730 11600 -22660
rect 11670 -22730 11710 -22660
rect 11780 -22730 11820 -22660
rect 11890 -22730 11930 -22660
rect 12000 -22730 12040 -22660
rect 12110 -22730 12150 -22660
rect 12220 -22730 12260 -22660
rect 12330 -22730 12370 -22660
rect 12440 -22730 12480 -22660
rect 12550 -22730 12590 -22660
rect 12660 -22730 12690 -22660
rect 11090 -22770 12690 -22730
rect 11090 -22840 11160 -22770
rect 11230 -22840 11270 -22770
rect 11340 -22840 11380 -22770
rect 11450 -22840 11490 -22770
rect 11560 -22840 11600 -22770
rect 11670 -22840 11710 -22770
rect 11780 -22840 11820 -22770
rect 11890 -22840 11930 -22770
rect 12000 -22840 12040 -22770
rect 12110 -22840 12150 -22770
rect 12220 -22840 12260 -22770
rect 12330 -22840 12370 -22770
rect 12440 -22840 12480 -22770
rect 12550 -22840 12590 -22770
rect 12660 -22840 12690 -22770
rect 11090 -22890 12690 -22840
<< via3 >>
rect -4730 8430 -4660 8500
rect -4640 8430 -4570 8500
rect -4550 8430 -4480 8500
rect -4460 8430 -4390 8500
rect -4370 8430 -4300 8500
rect -4280 8430 -4210 8500
rect -4190 8430 -4120 8500
rect -4100 8430 -4030 8500
rect -4010 8430 -3940 8500
rect -3920 8430 -3850 8500
rect -3830 8430 -3760 8500
rect -3740 8430 -3670 8500
rect -3650 8430 -3580 8500
rect -3560 8430 -3490 8500
rect -3470 8430 -3400 8500
rect -3380 8430 -3310 8500
rect -3290 8430 -3220 8500
rect -3200 8430 -3130 8500
rect -3110 8430 -3040 8500
rect -3020 8430 -2950 8500
rect -2930 8430 -2860 8500
rect -2840 8430 -2770 8500
rect -2750 8430 -2680 8500
rect -2660 8430 -2590 8500
rect -2570 8430 -2500 8500
rect -2480 8430 -2410 8500
rect -2390 8430 -2320 8500
rect -2300 8430 -2230 8500
rect -2210 8430 -2140 8500
rect -2120 8430 -2050 8500
rect -2030 8430 -1960 8500
rect -1940 8430 -1870 8500
rect -1850 8430 -1780 8500
rect -1720 8430 -1650 8500
rect -1630 8430 -1560 8500
rect -1540 8430 -1470 8500
rect -1450 8430 -1380 8500
rect -1360 8430 -1290 8500
rect -1270 8430 -1200 8500
rect -1180 8430 -1110 8500
rect -1090 8430 -1020 8500
rect -1000 8430 -930 8500
rect -910 8430 -840 8500
rect -820 8430 -750 8500
rect -730 8430 -660 8500
rect -640 8430 -570 8500
rect -550 8430 -480 8500
rect -460 8430 -390 8500
rect -370 8430 -300 8500
rect -280 8430 -210 8500
rect -190 8430 -120 8500
rect -100 8430 -30 8500
rect -10 8430 60 8500
rect 80 8430 150 8500
rect 170 8430 240 8500
rect 260 8430 330 8500
rect 350 8430 420 8500
rect 440 8430 510 8500
rect 530 8430 600 8500
rect 620 8430 690 8500
rect 710 8430 780 8500
rect 800 8430 870 8500
rect 890 8430 960 8500
rect 980 8430 1050 8500
rect 1070 8430 1140 8500
rect 1160 8430 1230 8500
rect 1290 8430 1360 8500
rect 1380 8430 1450 8500
rect 1470 8430 1540 8500
rect 1560 8430 1630 8500
rect 1650 8430 1720 8500
rect 1740 8430 1810 8500
rect 1830 8430 1900 8500
rect 1920 8430 1990 8500
rect 2010 8430 2080 8500
rect 2100 8430 2170 8500
rect 2190 8430 2260 8500
rect 2280 8430 2350 8500
rect 2370 8430 2440 8500
rect 2460 8430 2530 8500
rect 2550 8430 2620 8500
rect 2640 8430 2710 8500
rect 2730 8430 2800 8500
rect 2820 8430 2890 8500
rect 2910 8430 2980 8500
rect 3000 8430 3070 8500
rect 3090 8430 3160 8500
rect 3180 8430 3250 8500
rect 3270 8430 3340 8500
rect 3360 8430 3430 8500
rect 3450 8430 3520 8500
rect 3540 8430 3610 8500
rect 3630 8430 3700 8500
rect 3720 8430 3790 8500
rect 3810 8430 3880 8500
rect 3900 8430 3970 8500
rect 3990 8430 4060 8500
rect 4080 8430 4150 8500
rect 4170 8430 4240 8500
rect 4300 8430 4370 8500
rect 4390 8430 4460 8500
rect 4480 8430 4550 8500
rect 4570 8430 4640 8500
rect 4660 8430 4730 8500
rect 4750 8430 4820 8500
rect 4840 8430 4910 8500
rect 4930 8430 5000 8500
rect 5020 8430 5090 8500
rect 5110 8430 5180 8500
rect 5200 8430 5270 8500
rect 5290 8430 5360 8500
rect 5380 8430 5450 8500
rect 5470 8430 5540 8500
rect 5560 8430 5630 8500
rect 5650 8430 5720 8500
rect 5740 8430 5810 8500
rect 5830 8430 5900 8500
rect 5920 8430 5990 8500
rect 6010 8430 6080 8500
rect 6100 8430 6170 8500
rect 6190 8430 6260 8500
rect 6280 8430 6350 8500
rect 6370 8430 6440 8500
rect 6460 8430 6530 8500
rect 6550 8430 6620 8500
rect 6640 8430 6710 8500
rect 6730 8430 6800 8500
rect 6820 8430 6890 8500
rect 6910 8430 6980 8500
rect 7000 8430 7070 8500
rect 7090 8430 7160 8500
rect 7180 8430 7250 8500
rect -4730 8340 -4660 8410
rect -4640 8340 -4570 8410
rect -4550 8340 -4480 8410
rect -4460 8340 -4390 8410
rect -4370 8340 -4300 8410
rect -4280 8340 -4210 8410
rect -4190 8340 -4120 8410
rect -4100 8340 -4030 8410
rect -4010 8340 -3940 8410
rect -3920 8340 -3850 8410
rect -3830 8340 -3760 8410
rect -3740 8340 -3670 8410
rect -3650 8340 -3580 8410
rect -3560 8340 -3490 8410
rect -3470 8340 -3400 8410
rect -3380 8340 -3310 8410
rect -3290 8340 -3220 8410
rect -3200 8340 -3130 8410
rect -3110 8340 -3040 8410
rect -3020 8340 -2950 8410
rect -2930 8340 -2860 8410
rect -2840 8340 -2770 8410
rect -2750 8340 -2680 8410
rect -2660 8340 -2590 8410
rect -2570 8340 -2500 8410
rect -2480 8340 -2410 8410
rect -2390 8340 -2320 8410
rect -2300 8340 -2230 8410
rect -2210 8340 -2140 8410
rect -2120 8340 -2050 8410
rect -2030 8340 -1960 8410
rect -1940 8340 -1870 8410
rect -1850 8340 -1780 8410
rect -1720 8340 -1650 8410
rect -1630 8340 -1560 8410
rect -1540 8340 -1470 8410
rect -1450 8340 -1380 8410
rect -1360 8340 -1290 8410
rect -1270 8340 -1200 8410
rect -1180 8340 -1110 8410
rect -1090 8340 -1020 8410
rect -1000 8340 -930 8410
rect -910 8340 -840 8410
rect -820 8340 -750 8410
rect -730 8340 -660 8410
rect -640 8340 -570 8410
rect -550 8340 -480 8410
rect -460 8340 -390 8410
rect -370 8340 -300 8410
rect -280 8340 -210 8410
rect -190 8340 -120 8410
rect -100 8340 -30 8410
rect -10 8340 60 8410
rect 80 8340 150 8410
rect 170 8340 240 8410
rect 260 8340 330 8410
rect 350 8340 420 8410
rect 440 8340 510 8410
rect 530 8340 600 8410
rect 620 8340 690 8410
rect 710 8340 780 8410
rect 800 8340 870 8410
rect 890 8340 960 8410
rect 980 8340 1050 8410
rect 1070 8340 1140 8410
rect 1160 8340 1230 8410
rect 1290 8340 1360 8410
rect 1380 8340 1450 8410
rect 1470 8340 1540 8410
rect 1560 8340 1630 8410
rect 1650 8340 1720 8410
rect 1740 8340 1810 8410
rect 1830 8340 1900 8410
rect 1920 8340 1990 8410
rect 2010 8340 2080 8410
rect 2100 8340 2170 8410
rect 2190 8340 2260 8410
rect 2280 8340 2350 8410
rect 2370 8340 2440 8410
rect 2460 8340 2530 8410
rect 2550 8340 2620 8410
rect 2640 8340 2710 8410
rect 2730 8340 2800 8410
rect 2820 8340 2890 8410
rect 2910 8340 2980 8410
rect 3000 8340 3070 8410
rect 3090 8340 3160 8410
rect 3180 8340 3250 8410
rect 3270 8340 3340 8410
rect 3360 8340 3430 8410
rect 3450 8340 3520 8410
rect 3540 8340 3610 8410
rect 3630 8340 3700 8410
rect 3720 8340 3790 8410
rect 3810 8340 3880 8410
rect 3900 8340 3970 8410
rect 3990 8340 4060 8410
rect 4080 8340 4150 8410
rect 4170 8340 4240 8410
rect 4300 8340 4370 8410
rect 4390 8340 4460 8410
rect 4480 8340 4550 8410
rect 4570 8340 4640 8410
rect 4660 8340 4730 8410
rect 4750 8340 4820 8410
rect 4840 8340 4910 8410
rect 4930 8340 5000 8410
rect 5020 8340 5090 8410
rect 5110 8340 5180 8410
rect 5200 8340 5270 8410
rect 5290 8340 5360 8410
rect 5380 8340 5450 8410
rect 5470 8340 5540 8410
rect 5560 8340 5630 8410
rect 5650 8340 5720 8410
rect 5740 8340 5810 8410
rect 5830 8340 5900 8410
rect 5920 8340 5990 8410
rect 6010 8340 6080 8410
rect 6100 8340 6170 8410
rect 6190 8340 6260 8410
rect 6280 8340 6350 8410
rect 6370 8340 6440 8410
rect 6460 8340 6530 8410
rect 6550 8340 6620 8410
rect 6640 8340 6710 8410
rect 6730 8340 6800 8410
rect 6820 8340 6890 8410
rect 6910 8340 6980 8410
rect 7000 8340 7070 8410
rect 7090 8340 7160 8410
rect 7180 8340 7250 8410
rect -4730 8250 -4660 8320
rect -4640 8250 -4570 8320
rect -4550 8250 -4480 8320
rect -4460 8250 -4390 8320
rect -4370 8250 -4300 8320
rect -4280 8250 -4210 8320
rect -4190 8250 -4120 8320
rect -4100 8250 -4030 8320
rect -4010 8250 -3940 8320
rect -3920 8250 -3850 8320
rect -3830 8250 -3760 8320
rect -3740 8250 -3670 8320
rect -3650 8250 -3580 8320
rect -3560 8250 -3490 8320
rect -3470 8250 -3400 8320
rect -3380 8250 -3310 8320
rect -3290 8250 -3220 8320
rect -3200 8250 -3130 8320
rect -3110 8250 -3040 8320
rect -3020 8250 -2950 8320
rect -2930 8250 -2860 8320
rect -2840 8250 -2770 8320
rect -2750 8250 -2680 8320
rect -2660 8250 -2590 8320
rect -2570 8250 -2500 8320
rect -2480 8250 -2410 8320
rect -2390 8250 -2320 8320
rect -2300 8250 -2230 8320
rect -2210 8250 -2140 8320
rect -2120 8250 -2050 8320
rect -2030 8250 -1960 8320
rect -1940 8250 -1870 8320
rect -1850 8250 -1780 8320
rect -1720 8250 -1650 8320
rect -1630 8250 -1560 8320
rect -1540 8250 -1470 8320
rect -1450 8250 -1380 8320
rect -1360 8250 -1290 8320
rect -1270 8250 -1200 8320
rect -1180 8250 -1110 8320
rect -1090 8250 -1020 8320
rect -1000 8250 -930 8320
rect -910 8250 -840 8320
rect -820 8250 -750 8320
rect -730 8250 -660 8320
rect -640 8250 -570 8320
rect -550 8250 -480 8320
rect -460 8250 -390 8320
rect -370 8250 -300 8320
rect -280 8250 -210 8320
rect -190 8250 -120 8320
rect -100 8250 -30 8320
rect -10 8250 60 8320
rect 80 8250 150 8320
rect 170 8250 240 8320
rect 260 8250 330 8320
rect 350 8250 420 8320
rect 440 8250 510 8320
rect 530 8250 600 8320
rect 620 8250 690 8320
rect 710 8250 780 8320
rect 800 8250 870 8320
rect 890 8250 960 8320
rect 980 8250 1050 8320
rect 1070 8250 1140 8320
rect 1160 8250 1230 8320
rect 1290 8250 1360 8320
rect 1380 8250 1450 8320
rect 1470 8250 1540 8320
rect 1560 8250 1630 8320
rect 1650 8250 1720 8320
rect 1740 8250 1810 8320
rect 1830 8250 1900 8320
rect 1920 8250 1990 8320
rect 2010 8250 2080 8320
rect 2100 8250 2170 8320
rect 2190 8250 2260 8320
rect 2280 8250 2350 8320
rect 2370 8250 2440 8320
rect 2460 8250 2530 8320
rect 2550 8250 2620 8320
rect 2640 8250 2710 8320
rect 2730 8250 2800 8320
rect 2820 8250 2890 8320
rect 2910 8250 2980 8320
rect 3000 8250 3070 8320
rect 3090 8250 3160 8320
rect 3180 8250 3250 8320
rect 3270 8250 3340 8320
rect 3360 8250 3430 8320
rect 3450 8250 3520 8320
rect 3540 8250 3610 8320
rect 3630 8250 3700 8320
rect 3720 8250 3790 8320
rect 3810 8250 3880 8320
rect 3900 8250 3970 8320
rect 3990 8250 4060 8320
rect 4080 8250 4150 8320
rect 4170 8250 4240 8320
rect 4300 8250 4370 8320
rect 4390 8250 4460 8320
rect 4480 8250 4550 8320
rect 4570 8250 4640 8320
rect 4660 8250 4730 8320
rect 4750 8250 4820 8320
rect 4840 8250 4910 8320
rect 4930 8250 5000 8320
rect 5020 8250 5090 8320
rect 5110 8250 5180 8320
rect 5200 8250 5270 8320
rect 5290 8250 5360 8320
rect 5380 8250 5450 8320
rect 5470 8250 5540 8320
rect 5560 8250 5630 8320
rect 5650 8250 5720 8320
rect 5740 8250 5810 8320
rect 5830 8250 5900 8320
rect 5920 8250 5990 8320
rect 6010 8250 6080 8320
rect 6100 8250 6170 8320
rect 6190 8250 6260 8320
rect 6280 8250 6350 8320
rect 6370 8250 6440 8320
rect 6460 8250 6530 8320
rect 6550 8250 6620 8320
rect 6640 8250 6710 8320
rect 6730 8250 6800 8320
rect 6820 8250 6890 8320
rect 6910 8250 6980 8320
rect 7000 8250 7070 8320
rect 7090 8250 7160 8320
rect 7180 8250 7250 8320
rect 7650 8430 7720 8500
rect 7740 8430 7810 8500
rect 7830 8430 7900 8500
rect 7920 8430 7990 8500
rect 8010 8430 8080 8500
rect 8100 8430 8170 8500
rect 8190 8430 8260 8500
rect 8280 8430 8350 8500
rect 8370 8430 8440 8500
rect 8460 8430 8530 8500
rect 8550 8430 8620 8500
rect 8640 8430 8710 8500
rect 8730 8430 8800 8500
rect 8820 8430 8890 8500
rect 8910 8430 8980 8500
rect 9000 8430 9070 8500
rect 9090 8430 9160 8500
rect 9180 8430 9250 8500
rect 9270 8430 9340 8500
rect 9360 8430 9430 8500
rect 9450 8430 9520 8500
rect 9540 8430 9610 8500
rect 9630 8430 9700 8500
rect 9720 8430 9790 8500
rect 9810 8430 9880 8500
rect 9900 8430 9970 8500
rect 9990 8430 10060 8500
rect 10080 8430 10150 8500
rect 10170 8430 10240 8500
rect 10260 8430 10330 8500
rect 10350 8430 10420 8500
rect 10440 8430 10510 8500
rect 10530 8430 10600 8500
rect 10660 8430 10730 8500
rect 10750 8430 10820 8500
rect 10840 8430 10910 8500
rect 10930 8430 11000 8500
rect 11020 8430 11090 8500
rect 11110 8430 11180 8500
rect 11200 8430 11270 8500
rect 11290 8430 11360 8500
rect 11380 8430 11450 8500
rect 11470 8430 11540 8500
rect 11560 8430 11630 8500
rect 11650 8430 11720 8500
rect 11740 8430 11810 8500
rect 11830 8430 11900 8500
rect 11920 8430 11990 8500
rect 12010 8430 12080 8500
rect 12100 8430 12170 8500
rect 12190 8430 12260 8500
rect 12280 8430 12350 8500
rect 12370 8430 12440 8500
rect 12460 8430 12530 8500
rect 12550 8430 12620 8500
rect 12640 8430 12710 8500
rect 12730 8430 12800 8500
rect 12820 8430 12890 8500
rect 12910 8430 12980 8500
rect 13000 8430 13070 8500
rect 13090 8430 13160 8500
rect 13180 8430 13250 8500
rect 13270 8430 13340 8500
rect 13360 8430 13430 8500
rect 13450 8430 13520 8500
rect 13540 8430 13610 8500
rect 13670 8430 13740 8500
rect 13760 8430 13830 8500
rect 13850 8430 13920 8500
rect 13940 8430 14010 8500
rect 14030 8430 14100 8500
rect 14120 8430 14190 8500
rect 14210 8430 14280 8500
rect 14300 8430 14370 8500
rect 14390 8430 14460 8500
rect 14480 8430 14550 8500
rect 14570 8430 14640 8500
rect 14660 8430 14730 8500
rect 14750 8430 14820 8500
rect 14840 8430 14910 8500
rect 14930 8430 15000 8500
rect 15020 8430 15090 8500
rect 15110 8430 15180 8500
rect 15200 8430 15270 8500
rect 15290 8430 15360 8500
rect 15380 8430 15450 8500
rect 15470 8430 15540 8500
rect 15560 8430 15630 8500
rect 15650 8430 15720 8500
rect 15740 8430 15810 8500
rect 15830 8430 15900 8500
rect 15920 8430 15990 8500
rect 16010 8430 16080 8500
rect 16100 8430 16170 8500
rect 16190 8430 16260 8500
rect 16280 8430 16350 8500
rect 16370 8430 16440 8500
rect 16460 8430 16530 8500
rect 16550 8430 16620 8500
rect 16680 8430 16750 8500
rect 16770 8430 16840 8500
rect 16860 8430 16930 8500
rect 16950 8430 17020 8500
rect 17040 8430 17110 8500
rect 17130 8430 17200 8500
rect 17220 8430 17290 8500
rect 17310 8430 17380 8500
rect 17400 8430 17470 8500
rect 17490 8430 17560 8500
rect 17580 8430 17650 8500
rect 17670 8430 17740 8500
rect 17760 8430 17830 8500
rect 17850 8430 17920 8500
rect 17940 8430 18010 8500
rect 18030 8430 18100 8500
rect 18120 8430 18190 8500
rect 18210 8430 18280 8500
rect 18300 8430 18370 8500
rect 18390 8430 18460 8500
rect 18480 8430 18550 8500
rect 18570 8430 18640 8500
rect 18660 8430 18730 8500
rect 18750 8430 18820 8500
rect 18840 8430 18910 8500
rect 18930 8430 19000 8500
rect 19020 8430 19090 8500
rect 19110 8430 19180 8500
rect 19200 8430 19270 8500
rect 19290 8430 19360 8500
rect 19380 8430 19450 8500
rect 19470 8430 19540 8500
rect 19560 8430 19630 8500
rect 7650 8340 7720 8410
rect 7740 8340 7810 8410
rect 7830 8340 7900 8410
rect 7920 8340 7990 8410
rect 8010 8340 8080 8410
rect 8100 8340 8170 8410
rect 8190 8340 8260 8410
rect 8280 8340 8350 8410
rect 8370 8340 8440 8410
rect 8460 8340 8530 8410
rect 8550 8340 8620 8410
rect 8640 8340 8710 8410
rect 8730 8340 8800 8410
rect 8820 8340 8890 8410
rect 8910 8340 8980 8410
rect 9000 8340 9070 8410
rect 9090 8340 9160 8410
rect 9180 8340 9250 8410
rect 9270 8340 9340 8410
rect 9360 8340 9430 8410
rect 9450 8340 9520 8410
rect 9540 8340 9610 8410
rect 9630 8340 9700 8410
rect 9720 8340 9790 8410
rect 9810 8340 9880 8410
rect 9900 8340 9970 8410
rect 9990 8340 10060 8410
rect 10080 8340 10150 8410
rect 10170 8340 10240 8410
rect 10260 8340 10330 8410
rect 10350 8340 10420 8410
rect 10440 8340 10510 8410
rect 10530 8340 10600 8410
rect 10660 8340 10730 8410
rect 10750 8340 10820 8410
rect 10840 8340 10910 8410
rect 10930 8340 11000 8410
rect 11020 8340 11090 8410
rect 11110 8340 11180 8410
rect 11200 8340 11270 8410
rect 11290 8340 11360 8410
rect 11380 8340 11450 8410
rect 11470 8340 11540 8410
rect 11560 8340 11630 8410
rect 11650 8340 11720 8410
rect 11740 8340 11810 8410
rect 11830 8340 11900 8410
rect 11920 8340 11990 8410
rect 12010 8340 12080 8410
rect 12100 8340 12170 8410
rect 12190 8340 12260 8410
rect 12280 8340 12350 8410
rect 12370 8340 12440 8410
rect 12460 8340 12530 8410
rect 12550 8340 12620 8410
rect 12640 8340 12710 8410
rect 12730 8340 12800 8410
rect 12820 8340 12890 8410
rect 12910 8340 12980 8410
rect 13000 8340 13070 8410
rect 13090 8340 13160 8410
rect 13180 8340 13250 8410
rect 13270 8340 13340 8410
rect 13360 8340 13430 8410
rect 13450 8340 13520 8410
rect 13540 8340 13610 8410
rect 13670 8340 13740 8410
rect 13760 8340 13830 8410
rect 13850 8340 13920 8410
rect 13940 8340 14010 8410
rect 14030 8340 14100 8410
rect 14120 8340 14190 8410
rect 14210 8340 14280 8410
rect 14300 8340 14370 8410
rect 14390 8340 14460 8410
rect 14480 8340 14550 8410
rect 14570 8340 14640 8410
rect 14660 8340 14730 8410
rect 14750 8340 14820 8410
rect 14840 8340 14910 8410
rect 14930 8340 15000 8410
rect 15020 8340 15090 8410
rect 15110 8340 15180 8410
rect 15200 8340 15270 8410
rect 15290 8340 15360 8410
rect 15380 8340 15450 8410
rect 15470 8340 15540 8410
rect 15560 8340 15630 8410
rect 15650 8340 15720 8410
rect 15740 8340 15810 8410
rect 15830 8340 15900 8410
rect 15920 8340 15990 8410
rect 16010 8340 16080 8410
rect 16100 8340 16170 8410
rect 16190 8340 16260 8410
rect 16280 8340 16350 8410
rect 16370 8340 16440 8410
rect 16460 8340 16530 8410
rect 16550 8340 16620 8410
rect 16680 8340 16750 8410
rect 16770 8340 16840 8410
rect 16860 8340 16930 8410
rect 16950 8340 17020 8410
rect 17040 8340 17110 8410
rect 17130 8340 17200 8410
rect 17220 8340 17290 8410
rect 17310 8340 17380 8410
rect 17400 8340 17470 8410
rect 17490 8340 17560 8410
rect 17580 8340 17650 8410
rect 17670 8340 17740 8410
rect 17760 8340 17830 8410
rect 17850 8340 17920 8410
rect 17940 8340 18010 8410
rect 18030 8340 18100 8410
rect 18120 8340 18190 8410
rect 18210 8340 18280 8410
rect 18300 8340 18370 8410
rect 18390 8340 18460 8410
rect 18480 8340 18550 8410
rect 18570 8340 18640 8410
rect 18660 8340 18730 8410
rect 18750 8340 18820 8410
rect 18840 8340 18910 8410
rect 18930 8340 19000 8410
rect 19020 8340 19090 8410
rect 19110 8340 19180 8410
rect 19200 8340 19270 8410
rect 19290 8340 19360 8410
rect 19380 8340 19450 8410
rect 19470 8340 19540 8410
rect 19560 8340 19630 8410
rect 7650 8250 7720 8320
rect 7740 8250 7810 8320
rect 7830 8250 7900 8320
rect 7920 8250 7990 8320
rect 8010 8250 8080 8320
rect 8100 8250 8170 8320
rect 8190 8250 8260 8320
rect 8280 8250 8350 8320
rect 8370 8250 8440 8320
rect 8460 8250 8530 8320
rect 8550 8250 8620 8320
rect 8640 8250 8710 8320
rect 8730 8250 8800 8320
rect 8820 8250 8890 8320
rect 8910 8250 8980 8320
rect 9000 8250 9070 8320
rect 9090 8250 9160 8320
rect 9180 8250 9250 8320
rect 9270 8250 9340 8320
rect 9360 8250 9430 8320
rect 9450 8250 9520 8320
rect 9540 8250 9610 8320
rect 9630 8250 9700 8320
rect 9720 8250 9790 8320
rect 9810 8250 9880 8320
rect 9900 8250 9970 8320
rect 9990 8250 10060 8320
rect 10080 8250 10150 8320
rect 10170 8250 10240 8320
rect 10260 8250 10330 8320
rect 10350 8250 10420 8320
rect 10440 8250 10510 8320
rect 10530 8250 10600 8320
rect 10660 8250 10730 8320
rect 10750 8250 10820 8320
rect 10840 8250 10910 8320
rect 10930 8250 11000 8320
rect 11020 8250 11090 8320
rect 11110 8250 11180 8320
rect 11200 8250 11270 8320
rect 11290 8250 11360 8320
rect 11380 8250 11450 8320
rect 11470 8250 11540 8320
rect 11560 8250 11630 8320
rect 11650 8250 11720 8320
rect 11740 8250 11810 8320
rect 11830 8250 11900 8320
rect 11920 8250 11990 8320
rect 12010 8250 12080 8320
rect 12100 8250 12170 8320
rect 12190 8250 12260 8320
rect 12280 8250 12350 8320
rect 12370 8250 12440 8320
rect 12460 8250 12530 8320
rect 12550 8250 12620 8320
rect 12640 8250 12710 8320
rect 12730 8250 12800 8320
rect 12820 8250 12890 8320
rect 12910 8250 12980 8320
rect 13000 8250 13070 8320
rect 13090 8250 13160 8320
rect 13180 8250 13250 8320
rect 13270 8250 13340 8320
rect 13360 8250 13430 8320
rect 13450 8250 13520 8320
rect 13540 8250 13610 8320
rect 13670 8250 13740 8320
rect 13760 8250 13830 8320
rect 13850 8250 13920 8320
rect 13940 8250 14010 8320
rect 14030 8250 14100 8320
rect 14120 8250 14190 8320
rect 14210 8250 14280 8320
rect 14300 8250 14370 8320
rect 14390 8250 14460 8320
rect 14480 8250 14550 8320
rect 14570 8250 14640 8320
rect 14660 8250 14730 8320
rect 14750 8250 14820 8320
rect 14840 8250 14910 8320
rect 14930 8250 15000 8320
rect 15020 8250 15090 8320
rect 15110 8250 15180 8320
rect 15200 8250 15270 8320
rect 15290 8250 15360 8320
rect 15380 8250 15450 8320
rect 15470 8250 15540 8320
rect 15560 8250 15630 8320
rect 15650 8250 15720 8320
rect 15740 8250 15810 8320
rect 15830 8250 15900 8320
rect 15920 8250 15990 8320
rect 16010 8250 16080 8320
rect 16100 8250 16170 8320
rect 16190 8250 16260 8320
rect 16280 8250 16350 8320
rect 16370 8250 16440 8320
rect 16460 8250 16530 8320
rect 16550 8250 16620 8320
rect 16680 8250 16750 8320
rect 16770 8250 16840 8320
rect 16860 8250 16930 8320
rect 16950 8250 17020 8320
rect 17040 8250 17110 8320
rect 17130 8250 17200 8320
rect 17220 8250 17290 8320
rect 17310 8250 17380 8320
rect 17400 8250 17470 8320
rect 17490 8250 17560 8320
rect 17580 8250 17650 8320
rect 17670 8250 17740 8320
rect 17760 8250 17830 8320
rect 17850 8250 17920 8320
rect 17940 8250 18010 8320
rect 18030 8250 18100 8320
rect 18120 8250 18190 8320
rect 18210 8250 18280 8320
rect 18300 8250 18370 8320
rect 18390 8250 18460 8320
rect 18480 8250 18550 8320
rect 18570 8250 18640 8320
rect 18660 8250 18730 8320
rect 18750 8250 18820 8320
rect 18840 8250 18910 8320
rect 18930 8250 19000 8320
rect 19020 8250 19090 8320
rect 19110 8250 19180 8320
rect 19200 8250 19270 8320
rect 19290 8250 19360 8320
rect 19380 8250 19450 8320
rect 19470 8250 19540 8320
rect 19560 8250 19630 8320
rect 7040 7840 7110 7910
rect 7140 7840 7210 7910
rect 7240 7840 7310 7910
rect 7040 7750 7110 7820
rect 7140 7750 7210 7820
rect 7240 7750 7310 7820
rect 1570 6780 1640 6850
rect 1680 6780 1750 6850
rect 1790 6780 1860 6850
rect 1900 6780 1970 6850
rect 2010 6780 2080 6850
rect 2120 6780 2190 6850
rect 2230 6780 2300 6850
rect 2340 6780 2410 6850
rect 2450 6780 2520 6850
rect 2560 6780 2630 6850
rect 2670 6780 2740 6850
rect 2780 6780 2850 6850
rect 2890 6780 2960 6850
rect 3000 6780 3070 6850
rect 1570 6670 1640 6740
rect 1680 6670 1750 6740
rect 1790 6670 1860 6740
rect 1900 6670 1970 6740
rect 2010 6670 2080 6740
rect 2120 6670 2190 6740
rect 2230 6670 2300 6740
rect 2340 6670 2410 6740
rect 2450 6670 2520 6740
rect 2560 6670 2630 6740
rect 2670 6670 2740 6740
rect 2780 6670 2850 6740
rect 2890 6670 2960 6740
rect 3000 6670 3070 6740
rect 7590 7840 7660 7910
rect 7690 7840 7760 7910
rect 7790 7840 7860 7910
rect 7590 7750 7660 7820
rect 7690 7750 7760 7820
rect 7790 7750 7860 7820
rect 7410 5320 7480 5390
rect 7410 5210 7480 5280
rect 7410 5100 7480 5170
rect 7410 4990 7480 5060
rect 7410 4880 7480 4950
rect 35790 7750 35860 7820
rect 35880 7750 35950 7820
rect 35970 7750 36040 7820
rect 35790 7660 35860 7730
rect 35880 7660 35950 7730
rect 35970 7660 36040 7730
rect 35790 7570 35860 7640
rect 35880 7570 35950 7640
rect 35970 7570 36040 7640
rect 35790 7480 35860 7550
rect 35880 7480 35950 7550
rect 35970 7480 36040 7550
rect 35790 7390 35860 7460
rect 35880 7390 35950 7460
rect 35970 7390 36040 7460
rect 35790 7300 35860 7370
rect 35880 7300 35950 7370
rect 35970 7300 36040 7370
rect 21090 7140 21160 7210
rect 21200 7140 21270 7210
rect 21310 7140 21380 7210
rect 21420 7140 21490 7210
rect 21090 7030 21160 7100
rect 21200 7030 21270 7100
rect 21310 7030 21380 7100
rect 21420 7030 21490 7100
rect 23490 7140 23560 7210
rect 23600 7140 23670 7210
rect 23710 7140 23780 7210
rect 23820 7140 23890 7210
rect 23490 7030 23560 7100
rect 23600 7030 23670 7100
rect 23710 7030 23780 7100
rect 23820 7030 23890 7100
rect 35790 7210 35860 7280
rect 35880 7210 35950 7280
rect 35970 7210 36040 7280
rect 35790 7080 35860 7150
rect 35880 7080 35950 7150
rect 35970 7080 36040 7150
rect 35790 6990 35860 7060
rect 35880 6990 35950 7060
rect 35970 6990 36040 7060
rect 11790 6810 11860 6880
rect 11900 6810 11970 6880
rect 12010 6810 12080 6880
rect 12120 6810 12190 6880
rect 12230 6810 12300 6880
rect 12340 6810 12410 6880
rect 12450 6810 12520 6880
rect 12560 6810 12630 6880
rect 12670 6810 12740 6880
rect 12780 6810 12850 6880
rect 12890 6810 12960 6880
rect 13000 6810 13070 6880
rect 13110 6810 13180 6880
rect 13220 6810 13290 6880
rect 11790 6700 11860 6770
rect 11900 6700 11970 6770
rect 12010 6700 12080 6770
rect 12120 6700 12190 6770
rect 12230 6700 12300 6770
rect 12340 6700 12410 6770
rect 12450 6700 12520 6770
rect 12560 6700 12630 6770
rect 12670 6700 12740 6770
rect 12780 6700 12850 6770
rect 12890 6700 12960 6770
rect 13000 6700 13070 6770
rect 13110 6700 13180 6770
rect 13220 6700 13290 6770
rect 35790 6900 35860 6970
rect 35880 6900 35950 6970
rect 35970 6900 36040 6970
rect 35790 6810 35860 6880
rect 35880 6810 35950 6880
rect 35970 6810 36040 6880
rect 35790 6720 35860 6790
rect 35880 6720 35950 6790
rect 35970 6720 36040 6790
rect 35790 6630 35860 6700
rect 35880 6630 35950 6700
rect 35970 6630 36040 6700
rect 35790 6540 35860 6610
rect 35880 6540 35950 6610
rect 35970 6540 36040 6610
rect 35790 6450 35860 6520
rect 35880 6450 35950 6520
rect 35970 6450 36040 6520
rect 35790 6360 35860 6430
rect 35880 6360 35950 6430
rect 35970 6360 36040 6430
rect 28340 6230 28410 6300
rect 28450 6230 28520 6300
rect 28340 6100 28410 6170
rect 28450 6100 28520 6170
rect 28340 5970 28410 6040
rect 28450 5970 28520 6040
rect 35790 6270 35860 6340
rect 35880 6270 35950 6340
rect 35970 6270 36040 6340
rect 35790 6180 35860 6250
rect 35880 6180 35950 6250
rect 35970 6180 36040 6250
rect 35790 6090 35860 6160
rect 35880 6090 35950 6160
rect 35970 6090 36040 6160
rect 35790 6000 35860 6070
rect 35880 6000 35950 6070
rect 35970 6000 36040 6070
rect 35790 5910 35860 5980
rect 35880 5910 35950 5980
rect 35970 5910 36040 5980
rect 35790 5820 35860 5890
rect 35880 5820 35950 5890
rect 35970 5820 36040 5890
rect 35790 5730 35860 5800
rect 35880 5730 35950 5800
rect 35970 5730 36040 5800
rect 35790 5640 35860 5710
rect 35880 5640 35950 5710
rect 35970 5640 36040 5710
rect 35790 5550 35860 5620
rect 35880 5550 35950 5620
rect 35970 5550 36040 5620
rect 35790 5460 35860 5530
rect 35880 5460 35950 5530
rect 35970 5460 36040 5530
rect 35790 5370 35860 5440
rect 35880 5370 35950 5440
rect 35970 5370 36040 5440
rect 35790 5280 35860 5350
rect 35880 5280 35950 5350
rect 35970 5280 36040 5350
rect 35790 5190 35860 5260
rect 35880 5190 35950 5260
rect 35970 5190 36040 5260
rect 35790 5100 35860 5170
rect 35880 5100 35950 5170
rect 35970 5100 36040 5170
rect 35790 5010 35860 5080
rect 35880 5010 35950 5080
rect 35970 5010 36040 5080
rect 35790 4920 35860 4990
rect 35880 4920 35950 4990
rect 35970 4920 36040 4990
rect 35790 4830 35860 4900
rect 35880 4830 35950 4900
rect 35970 4830 36040 4900
rect 35790 4740 35860 4810
rect 35880 4740 35950 4810
rect 35970 4740 36040 4810
rect 35790 4650 35860 4720
rect 35880 4650 35950 4720
rect 35970 4650 36040 4720
rect 35790 4560 35860 4630
rect 35880 4560 35950 4630
rect 35970 4560 36040 4630
rect 35790 4470 35860 4540
rect 35880 4470 35950 4540
rect 35970 4470 36040 4540
rect 35790 4380 35860 4450
rect 35880 4380 35950 4450
rect 35970 4380 36040 4450
rect 35790 4290 35860 4360
rect 35880 4290 35950 4360
rect 35970 4290 36040 4360
rect 35790 4200 35860 4270
rect 35880 4200 35950 4270
rect 35970 4200 36040 4270
rect 35790 4070 35860 4140
rect 35880 4070 35950 4140
rect 35970 4070 36040 4140
rect 35790 3980 35860 4050
rect 35880 3980 35950 4050
rect 35970 3980 36040 4050
rect 35790 3890 35860 3960
rect 35880 3890 35950 3960
rect 35970 3890 36040 3960
rect 35790 3800 35860 3870
rect 35880 3800 35950 3870
rect 35970 3800 36040 3870
rect 35790 3710 35860 3780
rect 35880 3710 35950 3780
rect 35970 3710 36040 3780
rect 35790 3620 35860 3690
rect 35880 3620 35950 3690
rect 35970 3620 36040 3690
rect 35790 3530 35860 3600
rect 35880 3530 35950 3600
rect 35970 3530 36040 3600
rect 35790 3440 35860 3510
rect 35880 3440 35950 3510
rect 35970 3440 36040 3510
rect 22320 3290 22390 3360
rect 22430 3290 22500 3360
rect 22540 3290 22610 3360
rect 22320 3180 22390 3250
rect 22430 3180 22500 3250
rect 22540 3180 22610 3250
rect 22320 3070 22390 3140
rect 22430 3070 22500 3140
rect 22540 3070 22610 3140
rect 35790 3350 35860 3420
rect 35880 3350 35950 3420
rect 35970 3350 36040 3420
rect 35790 3260 35860 3330
rect 35880 3260 35950 3330
rect 35970 3260 36040 3330
rect 35790 3170 35860 3240
rect 35880 3170 35950 3240
rect 35970 3170 36040 3240
rect 35790 3080 35860 3150
rect 35880 3080 35950 3150
rect 35970 3080 36040 3150
rect 35790 2990 35860 3060
rect 35880 2990 35950 3060
rect 35970 2990 36040 3060
rect 1150 -860 1220 -790
rect 1260 -860 1330 -790
rect 1370 -860 1440 -790
rect 1480 -860 1550 -790
rect 1590 -860 1660 -790
rect 1700 -860 1770 -790
rect 1810 -860 1880 -790
rect 1920 -860 1990 -790
rect 2030 -860 2100 -790
rect 2140 -860 2210 -790
rect 2250 -860 2320 -790
rect 2360 -860 2430 -790
rect 2470 -860 2540 -790
rect 2580 -860 2650 -790
rect 1150 -970 1220 -900
rect 1260 -970 1330 -900
rect 1370 -970 1440 -900
rect 1480 -970 1550 -900
rect 1590 -970 1660 -900
rect 1700 -970 1770 -900
rect 1810 -970 1880 -900
rect 1920 -970 1990 -900
rect 2030 -970 2100 -900
rect 2140 -970 2210 -900
rect 2250 -970 2320 -900
rect 2360 -970 2430 -900
rect 2470 -970 2540 -900
rect 2580 -970 2650 -900
rect 1570 -2850 1640 -2780
rect 1680 -2850 1750 -2780
rect 1790 -2850 1860 -2780
rect 1900 -2850 1970 -2780
rect 2010 -2850 2080 -2780
rect 2120 -2850 2190 -2780
rect 2230 -2850 2300 -2780
rect 2340 -2850 2410 -2780
rect 2450 -2850 2520 -2780
rect 2560 -2850 2630 -2780
rect 2670 -2850 2740 -2780
rect 2780 -2850 2850 -2780
rect 2890 -2850 2960 -2780
rect 3000 -2850 3070 -2780
rect 1570 -2960 1640 -2890
rect 1680 -2960 1750 -2890
rect 1790 -2960 1860 -2890
rect 1900 -2960 1970 -2890
rect 2010 -2960 2080 -2890
rect 2120 -2960 2190 -2890
rect 2230 -2960 2300 -2890
rect 2340 -2960 2410 -2890
rect 2450 -2960 2520 -2890
rect 2560 -2960 2630 -2890
rect 2670 -2960 2740 -2890
rect 2780 -2960 2850 -2890
rect 2890 -2960 2960 -2890
rect 3000 -2960 3070 -2890
rect -160 -4300 -90 -4230
rect -70 -4300 0 -4230
rect 20 -4300 90 -4230
rect -160 -4390 -90 -4320
rect -70 -4390 0 -4320
rect 20 -4390 90 -4320
rect -160 -4480 -90 -4410
rect -70 -4480 0 -4410
rect 20 -4480 90 -4410
rect -160 -4570 -90 -4500
rect -70 -4570 0 -4500
rect 20 -4570 90 -4500
rect -160 -4660 -90 -4590
rect -70 -4660 0 -4590
rect 20 -4660 90 -4590
rect -160 -4750 -90 -4680
rect -70 -4750 0 -4680
rect 20 -4750 90 -4680
rect -160 -4840 -90 -4770
rect -70 -4840 0 -4770
rect 20 -4840 90 -4770
rect -160 -4930 -90 -4860
rect -70 -4930 0 -4860
rect 20 -4930 90 -4860
rect -160 -5020 -90 -4950
rect -70 -5020 0 -4950
rect 20 -5020 90 -4950
rect -160 -5110 -90 -5040
rect -70 -5110 0 -5040
rect 20 -5110 90 -5040
rect -160 -5200 -90 -5130
rect -70 -5200 0 -5130
rect 20 -5200 90 -5130
rect -2140 -5310 -2070 -5240
rect -2030 -5310 -1960 -5240
rect -2140 -5420 -2070 -5350
rect -2030 -5420 -1960 -5350
rect -2140 -5530 -2070 -5460
rect -2030 -5530 -1960 -5460
rect -2140 -5640 -2070 -5570
rect -2030 -5640 -1960 -5570
rect -160 -5290 -90 -5220
rect -70 -5290 0 -5220
rect 20 -5290 90 -5220
rect -160 -5380 -90 -5310
rect -70 -5380 0 -5310
rect 20 -5380 90 -5310
rect -160 -5470 -90 -5400
rect -70 -5470 0 -5400
rect 20 -5470 90 -5400
rect 35790 2900 35860 2970
rect 35880 2900 35950 2970
rect 35970 2900 36040 2970
rect 35790 2810 35860 2880
rect 35880 2810 35950 2880
rect 35970 2810 36040 2880
rect 35790 2720 35860 2790
rect 35880 2720 35950 2790
rect 35970 2720 36040 2790
rect 35790 2630 35860 2700
rect 35880 2630 35950 2700
rect 35970 2630 36040 2700
rect 20070 2530 20140 2600
rect 20180 2530 20250 2600
rect 20290 2530 20360 2600
rect 20400 2530 20470 2600
rect 20070 2420 20140 2490
rect 20180 2420 20250 2490
rect 20290 2420 20360 2490
rect 20400 2420 20470 2490
rect 24550 2530 24620 2600
rect 24660 2530 24730 2600
rect 24770 2530 24840 2600
rect 24880 2530 24950 2600
rect 24550 2420 24620 2490
rect 24660 2420 24730 2490
rect 24770 2420 24840 2490
rect 24880 2420 24950 2490
rect 35790 2540 35860 2610
rect 35880 2540 35950 2610
rect 35970 2540 36040 2610
rect 35790 2450 35860 2520
rect 35880 2450 35950 2520
rect 35970 2450 36040 2520
rect 35790 2360 35860 2430
rect 35880 2360 35950 2430
rect 35970 2360 36040 2430
rect 35790 2270 35860 2340
rect 35880 2270 35950 2340
rect 35970 2270 36040 2340
rect 35790 2180 35860 2250
rect 35880 2180 35950 2250
rect 35970 2180 36040 2250
rect 35790 2090 35860 2160
rect 35880 2090 35950 2160
rect 35970 2090 36040 2160
rect 35790 2000 35860 2070
rect 35880 2000 35950 2070
rect 35970 2000 36040 2070
rect 35790 1910 35860 1980
rect 35880 1910 35950 1980
rect 35970 1910 36040 1980
rect 35790 1820 35860 1890
rect 35880 1820 35950 1890
rect 35970 1820 36040 1890
rect 35790 1730 35860 1800
rect 35880 1730 35950 1800
rect 35970 1730 36040 1800
rect 35790 1640 35860 1710
rect 35880 1640 35950 1710
rect 35970 1640 36040 1710
rect 35790 1550 35860 1620
rect 35880 1550 35950 1620
rect 35970 1550 36040 1620
rect 35790 1460 35860 1530
rect 35880 1460 35950 1530
rect 35970 1460 36040 1530
rect 35790 1370 35860 1440
rect 35880 1370 35950 1440
rect 35970 1370 36040 1440
rect 35790 1280 35860 1350
rect 35880 1280 35950 1350
rect 35970 1280 36040 1350
rect 35790 1190 35860 1260
rect 35880 1190 35950 1260
rect 35970 1190 36040 1260
rect 14600 1090 14670 1160
rect 14700 1090 14770 1160
rect 14810 1090 14880 1160
rect 14600 980 14670 1050
rect 14700 980 14770 1050
rect 14810 980 14880 1050
rect 14600 870 14670 940
rect 14700 870 14770 940
rect 14810 870 14880 940
rect 21090 850 21160 920
rect 21200 850 21270 920
rect 21310 850 21380 920
rect 21420 850 21490 920
rect 21090 740 21160 810
rect 21200 740 21270 810
rect 21310 740 21380 810
rect 21420 740 21490 810
rect 23490 850 23560 920
rect 23600 850 23670 920
rect 23710 850 23780 920
rect 23820 850 23890 920
rect 23490 740 23560 810
rect 23600 740 23670 810
rect 23710 740 23780 810
rect 23820 740 23890 810
rect 35790 150 35860 220
rect 35880 150 35950 220
rect 35970 150 36040 220
rect 35790 60 35860 130
rect 35880 60 35950 130
rect 35970 60 36040 130
rect 28340 -70 28410 0
rect 28450 -70 28520 0
rect 28340 -200 28410 -130
rect 28450 -200 28520 -130
rect 28340 -330 28410 -260
rect 28450 -330 28520 -260
rect 35790 -30 35860 40
rect 35880 -30 35950 40
rect 35970 -30 36040 40
rect 35790 -120 35860 -50
rect 35880 -120 35950 -50
rect 35970 -120 36040 -50
rect 35790 -210 35860 -140
rect 35880 -210 35950 -140
rect 35970 -210 36040 -140
rect 35790 -300 35860 -230
rect 35880 -300 35950 -230
rect 35970 -300 36040 -230
rect 7310 -4630 7380 -4560
rect 7420 -4630 7490 -4560
rect 7530 -4630 7600 -4560
rect 7310 -4740 7380 -4670
rect 7420 -4740 7490 -4670
rect 7530 -4740 7600 -4670
rect 7310 -4850 7380 -4780
rect 7420 -4850 7490 -4780
rect 7530 -4850 7600 -4780
rect 35790 -390 35860 -320
rect 35880 -390 35950 -320
rect 35970 -390 36040 -320
rect 35790 -520 35860 -450
rect 35880 -520 35950 -450
rect 35970 -520 36040 -450
rect 35790 -610 35860 -540
rect 35880 -610 35950 -540
rect 35970 -610 36040 -540
rect 35790 -700 35860 -630
rect 35880 -700 35950 -630
rect 35970 -700 36040 -630
rect 12250 -860 12320 -790
rect 12360 -860 12430 -790
rect 12470 -860 12540 -790
rect 12580 -860 12650 -790
rect 12690 -860 12760 -790
rect 12800 -860 12870 -790
rect 12910 -860 12980 -790
rect 13020 -860 13090 -790
rect 13130 -860 13200 -790
rect 13240 -860 13310 -790
rect 13350 -860 13420 -790
rect 13460 -860 13530 -790
rect 13570 -860 13640 -790
rect 13680 -860 13750 -790
rect 12250 -970 12320 -900
rect 12360 -970 12430 -900
rect 12470 -970 12540 -900
rect 12580 -970 12650 -900
rect 12690 -970 12760 -900
rect 12800 -970 12870 -900
rect 12910 -970 12980 -900
rect 13020 -970 13090 -900
rect 13130 -970 13200 -900
rect 13240 -970 13310 -900
rect 13350 -970 13420 -900
rect 13460 -970 13530 -900
rect 13570 -970 13640 -900
rect 13680 -970 13750 -900
rect 35790 -790 35860 -720
rect 35880 -790 35950 -720
rect 35970 -790 36040 -720
rect 35790 -880 35860 -810
rect 35880 -880 35950 -810
rect 35970 -880 36040 -810
rect 35790 -970 35860 -900
rect 35880 -970 35950 -900
rect 35970 -970 36040 -900
rect 35790 -1060 35860 -990
rect 35880 -1060 35950 -990
rect 35970 -1060 36040 -990
rect 35790 -1150 35860 -1080
rect 35880 -1150 35950 -1080
rect 35970 -1150 36040 -1080
rect 35790 -1240 35860 -1170
rect 35880 -1240 35950 -1170
rect 35970 -1240 36040 -1170
rect 35790 -1330 35860 -1260
rect 35880 -1330 35950 -1260
rect 35970 -1330 36040 -1260
rect 35790 -1420 35860 -1350
rect 35880 -1420 35950 -1350
rect 35970 -1420 36040 -1350
rect 35790 -1510 35860 -1440
rect 35880 -1510 35950 -1440
rect 35970 -1510 36040 -1440
rect 35790 -1600 35860 -1530
rect 35880 -1600 35950 -1530
rect 35970 -1600 36040 -1530
rect 35790 -1690 35860 -1620
rect 35880 -1690 35950 -1620
rect 35970 -1690 36040 -1620
rect 35790 -1780 35860 -1710
rect 35880 -1780 35950 -1710
rect 35970 -1780 36040 -1710
rect 35790 -1870 35860 -1800
rect 35880 -1870 35950 -1800
rect 35970 -1870 36040 -1800
rect 35790 -1960 35860 -1890
rect 35880 -1960 35950 -1890
rect 35970 -1960 36040 -1890
rect 35790 -2050 35860 -1980
rect 35880 -2050 35950 -1980
rect 35970 -2050 36040 -1980
rect 35790 -2140 35860 -2070
rect 35880 -2140 35950 -2070
rect 35970 -2140 36040 -2070
rect 35790 -2230 35860 -2160
rect 35880 -2230 35950 -2160
rect 35970 -2230 36040 -2160
rect 35790 -2320 35860 -2250
rect 35880 -2320 35950 -2250
rect 35970 -2320 36040 -2250
rect 35790 -2410 35860 -2340
rect 35880 -2410 35950 -2340
rect 35970 -2410 36040 -2340
rect 35790 -2500 35860 -2430
rect 35880 -2500 35950 -2430
rect 35970 -2500 36040 -2430
rect 35790 -2590 35860 -2520
rect 35880 -2590 35950 -2520
rect 35970 -2590 36040 -2520
rect 35790 -2680 35860 -2610
rect 35880 -2680 35950 -2610
rect 35970 -2680 36040 -2610
rect 11790 -2850 11860 -2780
rect 11900 -2850 11970 -2780
rect 12010 -2850 12080 -2780
rect 12120 -2850 12190 -2780
rect 12230 -2850 12300 -2780
rect 12340 -2850 12410 -2780
rect 12450 -2850 12520 -2780
rect 12560 -2850 12630 -2780
rect 12670 -2850 12740 -2780
rect 12780 -2850 12850 -2780
rect 12890 -2850 12960 -2780
rect 13000 -2850 13070 -2780
rect 13110 -2850 13180 -2780
rect 13220 -2850 13290 -2780
rect 11790 -2960 11860 -2890
rect 11900 -2960 11970 -2890
rect 12010 -2960 12080 -2890
rect 12120 -2960 12190 -2890
rect 12230 -2960 12300 -2890
rect 12340 -2960 12410 -2890
rect 12450 -2960 12520 -2890
rect 12560 -2960 12630 -2890
rect 12670 -2960 12740 -2890
rect 12780 -2960 12850 -2890
rect 12890 -2960 12960 -2890
rect 13000 -2960 13070 -2890
rect 13110 -2960 13180 -2890
rect 13220 -2960 13290 -2890
rect 35790 -2770 35860 -2700
rect 35880 -2770 35950 -2700
rect 35970 -2770 36040 -2700
rect 35790 -2860 35860 -2790
rect 35880 -2860 35950 -2790
rect 35970 -2860 36040 -2790
rect 35790 -2950 35860 -2880
rect 35880 -2950 35950 -2880
rect 35970 -2950 36040 -2880
rect 22340 -3120 22410 -3050
rect 22450 -3120 22520 -3050
rect 22560 -3120 22630 -3050
rect 22340 -3230 22410 -3160
rect 22450 -3230 22520 -3160
rect 22560 -3230 22630 -3160
rect 22340 -3340 22410 -3270
rect 22450 -3340 22520 -3270
rect 22560 -3340 22630 -3270
rect 35790 -3040 35860 -2970
rect 35880 -3040 35950 -2970
rect 35970 -3040 36040 -2970
rect 35790 -3130 35860 -3060
rect 35880 -3130 35950 -3060
rect 35970 -3130 36040 -3060
rect 35790 -3220 35860 -3150
rect 35880 -3220 35950 -3150
rect 35970 -3220 36040 -3150
rect 35790 -3310 35860 -3240
rect 35880 -3310 35950 -3240
rect 35970 -3310 36040 -3240
rect 35790 -3400 35860 -3330
rect 35880 -3400 35950 -3330
rect 35970 -3400 36040 -3330
rect 35790 -3530 35860 -3460
rect 35880 -3530 35950 -3460
rect 35970 -3530 36040 -3460
rect 35790 -3620 35860 -3550
rect 35880 -3620 35950 -3550
rect 35970 -3620 36040 -3550
rect 20070 -3760 20140 -3690
rect 20180 -3760 20250 -3690
rect 20290 -3760 20360 -3690
rect 20400 -3760 20470 -3690
rect 20070 -3870 20140 -3800
rect 20180 -3870 20250 -3800
rect 20290 -3870 20360 -3800
rect 20400 -3870 20470 -3800
rect 24550 -3760 24620 -3690
rect 24660 -3760 24730 -3690
rect 24770 -3760 24840 -3690
rect 24880 -3760 24950 -3690
rect 24550 -3870 24620 -3800
rect 24660 -3870 24730 -3800
rect 24770 -3870 24840 -3800
rect 24880 -3870 24950 -3800
rect 35790 -3710 35860 -3640
rect 35880 -3710 35950 -3640
rect 35970 -3710 36040 -3640
rect 35790 -3800 35860 -3730
rect 35880 -3800 35950 -3730
rect 35970 -3800 36040 -3730
rect 35790 -3890 35860 -3820
rect 35880 -3890 35950 -3820
rect 35970 -3890 36040 -3820
rect 8200 -6220 8270 -6150
rect 8300 -6220 8370 -6150
rect 8400 -6220 8470 -6150
rect 8200 -6320 8270 -6250
rect 8300 -6320 8370 -6250
rect 8400 -6320 8470 -6250
rect 35790 -3980 35860 -3910
rect 35880 -3980 35950 -3910
rect 35970 -3980 36040 -3910
rect 35790 -4070 35860 -4000
rect 35880 -4070 35950 -4000
rect 35970 -4070 36040 -4000
rect 35790 -4160 35860 -4090
rect 35880 -4160 35950 -4090
rect 35970 -4160 36040 -4090
rect 35790 -4250 35860 -4180
rect 35880 -4250 35950 -4180
rect 35970 -4250 36040 -4180
rect 35790 -4340 35860 -4270
rect 35880 -4340 35950 -4270
rect 35970 -4340 36040 -4270
rect 35790 -4430 35860 -4360
rect 35880 -4430 35950 -4360
rect 35970 -4430 36040 -4360
rect 35790 -4520 35860 -4450
rect 35880 -4520 35950 -4450
rect 35970 -4520 36040 -4450
rect 35790 -4610 35860 -4540
rect 35880 -4610 35950 -4540
rect 35970 -4610 36040 -4540
rect 35790 -4700 35860 -4630
rect 35880 -4700 35950 -4630
rect 35970 -4700 36040 -4630
rect 35790 -4790 35860 -4720
rect 35880 -4790 35950 -4720
rect 35970 -4790 36040 -4720
rect 35790 -4880 35860 -4810
rect 35880 -4880 35950 -4810
rect 35970 -4880 36040 -4810
rect 35790 -4970 35860 -4900
rect 35880 -4970 35950 -4900
rect 35970 -4970 36040 -4900
rect 35790 -5060 35860 -4990
rect 35880 -5060 35950 -4990
rect 35970 -5060 36040 -4990
rect 35790 -5150 35860 -5080
rect 35880 -5150 35950 -5080
rect 35970 -5150 36040 -5080
rect 35790 -5240 35860 -5170
rect 35880 -5240 35950 -5170
rect 35970 -5240 36040 -5170
rect 35790 -5330 35860 -5260
rect 35880 -5330 35950 -5260
rect 35970 -5330 36040 -5260
rect 35790 -5420 35860 -5350
rect 35880 -5420 35950 -5350
rect 35970 -5420 36040 -5350
rect 35790 -5510 35860 -5440
rect 35880 -5510 35950 -5440
rect 35970 -5510 36040 -5440
rect 35790 -5600 35860 -5530
rect 35880 -5600 35950 -5530
rect 35970 -5600 36040 -5530
rect 35790 -5690 35860 -5620
rect 35880 -5690 35950 -5620
rect 35970 -5690 36040 -5620
rect 35790 -5780 35860 -5710
rect 35880 -5780 35950 -5710
rect 35970 -5780 36040 -5710
rect 35790 -5870 35860 -5800
rect 35880 -5870 35950 -5800
rect 35970 -5870 36040 -5800
rect 35790 -5960 35860 -5890
rect 35880 -5960 35950 -5890
rect 35970 -5960 36040 -5890
rect 35790 -6050 35860 -5980
rect 35880 -6050 35950 -5980
rect 35970 -6050 36040 -5980
rect 35790 -6140 35860 -6070
rect 35880 -6140 35950 -6070
rect 35970 -6140 36040 -6070
rect 35790 -6230 35860 -6160
rect 35880 -6230 35950 -6160
rect 35970 -6230 36040 -6160
rect 35790 -6320 35860 -6250
rect 35880 -6320 35950 -6250
rect 35970 -6320 36040 -6250
rect 35790 -6410 35860 -6340
rect 35880 -6410 35950 -6340
rect 35970 -6410 36040 -6340
rect -160 -7700 -90 -7630
rect -70 -7700 0 -7630
rect 20 -7700 90 -7630
rect -160 -7790 -90 -7720
rect -70 -7790 0 -7720
rect 20 -7790 90 -7720
rect -2200 -7940 -2130 -7870
rect -2090 -7940 -2020 -7870
rect -2200 -8050 -2130 -7980
rect -2090 -8050 -2020 -7980
rect -2200 -8160 -2130 -8090
rect -2090 -8160 -2020 -8090
rect -2200 -8270 -2130 -8200
rect -2090 -8270 -2020 -8200
rect -160 -7880 -90 -7810
rect -70 -7880 0 -7810
rect 20 -7880 90 -7810
rect -160 -7970 -90 -7900
rect -70 -7970 0 -7900
rect 20 -7970 90 -7900
rect -160 -8060 -90 -7990
rect -70 -8060 0 -7990
rect 20 -8060 90 -7990
rect -160 -8150 -90 -8080
rect -70 -8150 0 -8080
rect 20 -8150 90 -8080
rect -160 -8240 -90 -8170
rect -70 -8240 0 -8170
rect 20 -8240 90 -8170
rect -160 -8330 -90 -8260
rect -70 -8330 0 -8260
rect 20 -8330 90 -8260
rect -160 -8420 -90 -8350
rect -70 -8420 0 -8350
rect 20 -8420 90 -8350
rect -160 -8510 -90 -8440
rect -70 -8510 0 -8440
rect 20 -8510 90 -8440
rect -160 -8600 -90 -8530
rect -70 -8600 0 -8530
rect 20 -8600 90 -8530
rect -2140 -8710 -2070 -8640
rect -2030 -8710 -1960 -8640
rect -2140 -8820 -2070 -8750
rect -2030 -8820 -1960 -8750
rect -2140 -8930 -2070 -8860
rect -2030 -8930 -1960 -8860
rect -2140 -9040 -2070 -8970
rect -2030 -9040 -1960 -8970
rect -160 -8690 -90 -8620
rect -70 -8690 0 -8620
rect 20 -8690 90 -8620
rect -160 -8780 -90 -8710
rect -70 -8780 0 -8710
rect 20 -8780 90 -8710
rect -160 -8870 -90 -8800
rect -70 -8870 0 -8800
rect 20 -8870 90 -8800
rect 1150 -10410 1220 -10340
rect 1260 -10410 1330 -10340
rect 1370 -10410 1440 -10340
rect 1480 -10410 1550 -10340
rect 1590 -10410 1660 -10340
rect 1700 -10410 1770 -10340
rect 1810 -10410 1880 -10340
rect 1920 -10410 1990 -10340
rect 2030 -10410 2100 -10340
rect 2140 -10410 2210 -10340
rect 2250 -10410 2320 -10340
rect 2360 -10410 2430 -10340
rect 2470 -10410 2540 -10340
rect 2580 -10410 2650 -10340
rect 1150 -10520 1220 -10450
rect 1260 -10520 1330 -10450
rect 1370 -10520 1440 -10450
rect 1480 -10520 1550 -10450
rect 1590 -10520 1660 -10450
rect 1700 -10520 1770 -10450
rect 1810 -10520 1880 -10450
rect 1920 -10520 1990 -10450
rect 2030 -10520 2100 -10450
rect 2140 -10520 2210 -10450
rect 2250 -10520 2320 -10450
rect 2360 -10520 2430 -10450
rect 2470 -10520 2540 -10450
rect 2580 -10520 2650 -10450
rect 2240 -12370 2310 -12300
rect 2350 -12370 2420 -12300
rect 2460 -12370 2530 -12300
rect 2570 -12370 2640 -12300
rect 2680 -12370 2750 -12300
rect 2790 -12370 2860 -12300
rect 2900 -12370 2970 -12300
rect 3010 -12370 3080 -12300
rect 3120 -12370 3190 -12300
rect 3230 -12370 3300 -12300
rect 3340 -12370 3410 -12300
rect 3450 -12370 3520 -12300
rect 3560 -12370 3630 -12300
rect 3670 -12370 3740 -12300
rect 2240 -12480 2310 -12410
rect 2350 -12480 2420 -12410
rect 2460 -12480 2530 -12410
rect 2570 -12480 2640 -12410
rect 2680 -12480 2750 -12410
rect 2790 -12480 2860 -12410
rect 2900 -12480 2970 -12410
rect 3010 -12480 3080 -12410
rect 3120 -12480 3190 -12410
rect 3230 -12480 3300 -12410
rect 3340 -12480 3410 -12410
rect 3450 -12480 3520 -12410
rect 3560 -12480 3630 -12410
rect 3670 -12480 3740 -12410
rect 8730 -8320 8800 -8250
rect 8830 -8320 8900 -8250
rect 8930 -8320 9000 -8250
rect 8730 -8420 8800 -8350
rect 8830 -8420 8900 -8350
rect 8930 -8420 9000 -8350
rect 14600 -8300 14670 -8230
rect 14700 -8300 14770 -8230
rect 14810 -8300 14880 -8230
rect 14600 -8410 14670 -8340
rect 14700 -8410 14770 -8340
rect 14810 -8410 14880 -8340
rect 14600 -8520 14670 -8450
rect 14700 -8520 14770 -8450
rect 14810 -8520 14880 -8450
rect 19230 -8630 19300 -8560
rect 19330 -8630 19400 -8560
rect 19430 -8630 19500 -8560
rect 19230 -8730 19300 -8660
rect 19330 -8730 19400 -8660
rect 19430 -8730 19500 -8660
rect 19230 -8830 19300 -8760
rect 19330 -8830 19400 -8760
rect 19430 -8830 19500 -8760
rect 19960 -9070 20030 -9000
rect 20060 -9070 20130 -9000
rect 20160 -9070 20230 -9000
rect 19960 -9170 20030 -9100
rect 20060 -9170 20130 -9100
rect 20160 -9170 20230 -9100
rect 19960 -9270 20030 -9200
rect 20060 -9270 20130 -9200
rect 20160 -9270 20230 -9200
rect 12290 -10440 12360 -10370
rect 12400 -10440 12470 -10370
rect 12510 -10440 12580 -10370
rect 12620 -10440 12690 -10370
rect 12730 -10440 12800 -10370
rect 12840 -10440 12910 -10370
rect 12950 -10440 13020 -10370
rect 13060 -10440 13130 -10370
rect 13170 -10440 13240 -10370
rect 13280 -10440 13350 -10370
rect 13390 -10440 13460 -10370
rect 13500 -10440 13570 -10370
rect 13610 -10440 13680 -10370
rect 13720 -10440 13790 -10370
rect 12290 -10550 12360 -10480
rect 12400 -10550 12470 -10480
rect 12510 -10550 12580 -10480
rect 12620 -10550 12690 -10480
rect 12730 -10550 12800 -10480
rect 12840 -10550 12910 -10480
rect 12950 -10550 13020 -10480
rect 13060 -10550 13130 -10480
rect 13170 -10550 13240 -10480
rect 13280 -10550 13350 -10480
rect 13390 -10550 13460 -10480
rect 13500 -10550 13570 -10480
rect 13610 -10550 13680 -10480
rect 13720 -10550 13790 -10480
rect 11120 -12370 11190 -12300
rect 11230 -12370 11300 -12300
rect 11340 -12370 11410 -12300
rect 11450 -12370 11520 -12300
rect 11560 -12370 11630 -12300
rect 11670 -12370 11740 -12300
rect 11780 -12370 11850 -12300
rect 11890 -12370 11960 -12300
rect 12000 -12370 12070 -12300
rect 12110 -12370 12180 -12300
rect 12220 -12370 12290 -12300
rect 12330 -12370 12400 -12300
rect 12440 -12370 12510 -12300
rect 12550 -12370 12620 -12300
rect 11120 -12480 11190 -12410
rect 11230 -12480 11300 -12410
rect 11340 -12480 11410 -12410
rect 11450 -12480 11520 -12410
rect 11560 -12480 11630 -12410
rect 11670 -12480 11740 -12410
rect 11780 -12480 11850 -12410
rect 11890 -12480 11960 -12410
rect 12000 -12480 12070 -12410
rect 12110 -12480 12180 -12410
rect 12220 -12480 12290 -12410
rect 12330 -12480 12400 -12410
rect 12440 -12480 12510 -12410
rect 12550 -12480 12620 -12410
rect 19230 -14290 19300 -14220
rect 19330 -14290 19400 -14220
rect 19430 -14290 19500 -14220
rect 19230 -14390 19300 -14320
rect 19330 -14390 19400 -14320
rect 19430 -14390 19500 -14320
rect 19230 -14490 19300 -14420
rect 19330 -14490 19400 -14420
rect 19430 -14490 19500 -14420
rect 20480 -14940 20550 -14870
rect 20580 -14940 20650 -14870
rect 20680 -14940 20750 -14870
rect 20480 -15040 20550 -14970
rect 20580 -15040 20650 -14970
rect 20680 -15040 20750 -14970
rect 20480 -15140 20550 -15070
rect 20580 -15140 20650 -15070
rect 20680 -15140 20750 -15070
rect 2280 -22730 2350 -22660
rect 2390 -22730 2460 -22660
rect 2500 -22730 2570 -22660
rect 2610 -22730 2680 -22660
rect 2720 -22730 2790 -22660
rect 2830 -22730 2900 -22660
rect 2940 -22730 3010 -22660
rect 3050 -22730 3120 -22660
rect 3160 -22730 3230 -22660
rect 3270 -22730 3340 -22660
rect 3380 -22730 3450 -22660
rect 3490 -22730 3560 -22660
rect 3600 -22730 3670 -22660
rect 3710 -22730 3780 -22660
rect 2280 -22840 2350 -22770
rect 2390 -22840 2460 -22770
rect 2500 -22840 2570 -22770
rect 2610 -22840 2680 -22770
rect 2720 -22840 2790 -22770
rect 2830 -22840 2900 -22770
rect 2940 -22840 3010 -22770
rect 3050 -22840 3120 -22770
rect 3160 -22840 3230 -22770
rect 3270 -22840 3340 -22770
rect 3380 -22840 3450 -22770
rect 3490 -22840 3560 -22770
rect 3600 -22840 3670 -22770
rect 3710 -22840 3780 -22770
rect 7230 -17670 7300 -17600
rect 7340 -17670 7410 -17600
rect 7450 -17670 7520 -17600
rect 7560 -17670 7630 -17600
rect 7230 -17780 7300 -17710
rect 7340 -17780 7410 -17710
rect 7450 -17780 7520 -17710
rect 7560 -17780 7630 -17710
rect 7230 -17890 7300 -17820
rect 7340 -17890 7410 -17820
rect 7450 -17890 7520 -17820
rect 7560 -17890 7630 -17820
rect 7230 -18000 7300 -17930
rect 7340 -18000 7410 -17930
rect 7450 -18000 7520 -17930
rect 7560 -18000 7630 -17930
rect 19230 -20360 19300 -20290
rect 19330 -20360 19400 -20290
rect 19430 -20360 19500 -20290
rect 19230 -20460 19300 -20390
rect 19330 -20460 19400 -20390
rect 19430 -20460 19500 -20390
rect 19230 -20560 19300 -20490
rect 19330 -20560 19400 -20490
rect 19430 -20560 19500 -20490
rect 20040 -20790 20110 -20720
rect 20140 -20790 20210 -20720
rect 20240 -20790 20310 -20720
rect 20040 -20890 20110 -20820
rect 20140 -20890 20210 -20820
rect 20240 -20890 20310 -20820
rect 20040 -20990 20110 -20920
rect 20140 -20990 20210 -20920
rect 20240 -20990 20310 -20920
rect 11160 -22730 11230 -22660
rect 11270 -22730 11340 -22660
rect 11380 -22730 11450 -22660
rect 11490 -22730 11560 -22660
rect 11600 -22730 11670 -22660
rect 11710 -22730 11780 -22660
rect 11820 -22730 11890 -22660
rect 11930 -22730 12000 -22660
rect 12040 -22730 12110 -22660
rect 12150 -22730 12220 -22660
rect 12260 -22730 12330 -22660
rect 12370 -22730 12440 -22660
rect 12480 -22730 12550 -22660
rect 12590 -22730 12660 -22660
rect 11160 -22840 11230 -22770
rect 11270 -22840 11340 -22770
rect 11380 -22840 11450 -22770
rect 11490 -22840 11560 -22770
rect 11600 -22840 11670 -22770
rect 11710 -22840 11780 -22770
rect 11820 -22840 11890 -22770
rect 11930 -22840 12000 -22770
rect 12040 -22840 12110 -22770
rect 12150 -22840 12220 -22770
rect 12260 -22840 12330 -22770
rect 12370 -22840 12440 -22770
rect 12480 -22840 12550 -22770
rect 12590 -22840 12660 -22770
<< mimcap >>
rect -4980 20790 7260 21110
rect -4980 20550 -4670 20790
rect -4430 20550 -4340 20790
rect -4100 20550 -4010 20790
rect -3770 20550 -3680 20790
rect -3440 20550 -3350 20790
rect -3110 20550 -3020 20790
rect -2780 20550 -2690 20790
rect -2450 20550 -2360 20790
rect -2120 20550 -2030 20790
rect -1790 20550 -1700 20790
rect -1460 20550 -1370 20790
rect -1130 20550 -1040 20790
rect -800 20550 -710 20790
rect -470 20550 -380 20790
rect -140 20550 -50 20790
rect 190 20550 280 20790
rect 520 20550 610 20790
rect 850 20550 940 20790
rect 1180 20550 1270 20790
rect 1510 20550 1600 20790
rect 1840 20550 1930 20790
rect 2170 20550 2260 20790
rect 2500 20550 2590 20790
rect 2830 20550 2920 20790
rect 3160 20550 3250 20790
rect 3490 20550 3580 20790
rect 3820 20550 3910 20790
rect 4150 20550 4240 20790
rect 4480 20550 4570 20790
rect 4810 20550 4900 20790
rect 5140 20550 5230 20790
rect 5470 20550 5560 20790
rect 5800 20550 5890 20790
rect 6130 20550 6220 20790
rect 6460 20550 6550 20790
rect 6790 20550 6880 20790
rect 7120 20550 7260 20790
rect -4980 20460 7260 20550
rect -4980 20220 -4670 20460
rect -4430 20220 -4340 20460
rect -4100 20220 -4010 20460
rect -3770 20220 -3680 20460
rect -3440 20220 -3350 20460
rect -3110 20220 -3020 20460
rect -2780 20220 -2690 20460
rect -2450 20220 -2360 20460
rect -2120 20220 -2030 20460
rect -1790 20220 -1700 20460
rect -1460 20220 -1370 20460
rect -1130 20220 -1040 20460
rect -800 20220 -710 20460
rect -470 20220 -380 20460
rect -140 20220 -50 20460
rect 190 20220 280 20460
rect 520 20220 610 20460
rect 850 20220 940 20460
rect 1180 20220 1270 20460
rect 1510 20220 1600 20460
rect 1840 20220 1930 20460
rect 2170 20220 2260 20460
rect 2500 20220 2590 20460
rect 2830 20220 2920 20460
rect 3160 20220 3250 20460
rect 3490 20220 3580 20460
rect 3820 20220 3910 20460
rect 4150 20220 4240 20460
rect 4480 20220 4570 20460
rect 4810 20220 4900 20460
rect 5140 20220 5230 20460
rect 5470 20220 5560 20460
rect 5800 20220 5890 20460
rect 6130 20220 6220 20460
rect 6460 20220 6550 20460
rect 6790 20220 6880 20460
rect 7120 20220 7260 20460
rect -4980 20130 7260 20220
rect -4980 19890 -4670 20130
rect -4430 19890 -4340 20130
rect -4100 19890 -4010 20130
rect -3770 19890 -3680 20130
rect -3440 19890 -3350 20130
rect -3110 19890 -3020 20130
rect -2780 19890 -2690 20130
rect -2450 19890 -2360 20130
rect -2120 19890 -2030 20130
rect -1790 19890 -1700 20130
rect -1460 19890 -1370 20130
rect -1130 19890 -1040 20130
rect -800 19890 -710 20130
rect -470 19890 -380 20130
rect -140 19890 -50 20130
rect 190 19890 280 20130
rect 520 19890 610 20130
rect 850 19890 940 20130
rect 1180 19890 1270 20130
rect 1510 19890 1600 20130
rect 1840 19890 1930 20130
rect 2170 19890 2260 20130
rect 2500 19890 2590 20130
rect 2830 19890 2920 20130
rect 3160 19890 3250 20130
rect 3490 19890 3580 20130
rect 3820 19890 3910 20130
rect 4150 19890 4240 20130
rect 4480 19890 4570 20130
rect 4810 19890 4900 20130
rect 5140 19890 5230 20130
rect 5470 19890 5560 20130
rect 5800 19890 5890 20130
rect 6130 19890 6220 20130
rect 6460 19890 6550 20130
rect 6790 19890 6880 20130
rect 7120 19890 7260 20130
rect -4980 19800 7260 19890
rect -4980 19560 -4670 19800
rect -4430 19560 -4340 19800
rect -4100 19560 -4010 19800
rect -3770 19560 -3680 19800
rect -3440 19560 -3350 19800
rect -3110 19560 -3020 19800
rect -2780 19560 -2690 19800
rect -2450 19560 -2360 19800
rect -2120 19560 -2030 19800
rect -1790 19560 -1700 19800
rect -1460 19560 -1370 19800
rect -1130 19560 -1040 19800
rect -800 19560 -710 19800
rect -470 19560 -380 19800
rect -140 19560 -50 19800
rect 190 19560 280 19800
rect 520 19560 610 19800
rect 850 19560 940 19800
rect 1180 19560 1270 19800
rect 1510 19560 1600 19800
rect 1840 19560 1930 19800
rect 2170 19560 2260 19800
rect 2500 19560 2590 19800
rect 2830 19560 2920 19800
rect 3160 19560 3250 19800
rect 3490 19560 3580 19800
rect 3820 19560 3910 19800
rect 4150 19560 4240 19800
rect 4480 19560 4570 19800
rect 4810 19560 4900 19800
rect 5140 19560 5230 19800
rect 5470 19560 5560 19800
rect 5800 19560 5890 19800
rect 6130 19560 6220 19800
rect 6460 19560 6550 19800
rect 6790 19560 6880 19800
rect 7120 19560 7260 19800
rect -4980 19470 7260 19560
rect -4980 19230 -4670 19470
rect -4430 19230 -4340 19470
rect -4100 19230 -4010 19470
rect -3770 19230 -3680 19470
rect -3440 19230 -3350 19470
rect -3110 19230 -3020 19470
rect -2780 19230 -2690 19470
rect -2450 19230 -2360 19470
rect -2120 19230 -2030 19470
rect -1790 19230 -1700 19470
rect -1460 19230 -1370 19470
rect -1130 19230 -1040 19470
rect -800 19230 -710 19470
rect -470 19230 -380 19470
rect -140 19230 -50 19470
rect 190 19230 280 19470
rect 520 19230 610 19470
rect 850 19230 940 19470
rect 1180 19230 1270 19470
rect 1510 19230 1600 19470
rect 1840 19230 1930 19470
rect 2170 19230 2260 19470
rect 2500 19230 2590 19470
rect 2830 19230 2920 19470
rect 3160 19230 3250 19470
rect 3490 19230 3580 19470
rect 3820 19230 3910 19470
rect 4150 19230 4240 19470
rect 4480 19230 4570 19470
rect 4810 19230 4900 19470
rect 5140 19230 5230 19470
rect 5470 19230 5560 19470
rect 5800 19230 5890 19470
rect 6130 19230 6220 19470
rect 6460 19230 6550 19470
rect 6790 19230 6880 19470
rect 7120 19230 7260 19470
rect -4980 19140 7260 19230
rect -4980 18900 -4670 19140
rect -4430 18900 -4340 19140
rect -4100 18900 -4010 19140
rect -3770 18900 -3680 19140
rect -3440 18900 -3350 19140
rect -3110 18900 -3020 19140
rect -2780 18900 -2690 19140
rect -2450 18900 -2360 19140
rect -2120 18900 -2030 19140
rect -1790 18900 -1700 19140
rect -1460 18900 -1370 19140
rect -1130 18900 -1040 19140
rect -800 18900 -710 19140
rect -470 18900 -380 19140
rect -140 18900 -50 19140
rect 190 18900 280 19140
rect 520 18900 610 19140
rect 850 18900 940 19140
rect 1180 18900 1270 19140
rect 1510 18900 1600 19140
rect 1840 18900 1930 19140
rect 2170 18900 2260 19140
rect 2500 18900 2590 19140
rect 2830 18900 2920 19140
rect 3160 18900 3250 19140
rect 3490 18900 3580 19140
rect 3820 18900 3910 19140
rect 4150 18900 4240 19140
rect 4480 18900 4570 19140
rect 4810 18900 4900 19140
rect 5140 18900 5230 19140
rect 5470 18900 5560 19140
rect 5800 18900 5890 19140
rect 6130 18900 6220 19140
rect 6460 18900 6550 19140
rect 6790 18900 6880 19140
rect 7120 18900 7260 19140
rect -4980 18810 7260 18900
rect -4980 18570 -4670 18810
rect -4430 18570 -4340 18810
rect -4100 18570 -4010 18810
rect -3770 18570 -3680 18810
rect -3440 18570 -3350 18810
rect -3110 18570 -3020 18810
rect -2780 18570 -2690 18810
rect -2450 18570 -2360 18810
rect -2120 18570 -2030 18810
rect -1790 18570 -1700 18810
rect -1460 18570 -1370 18810
rect -1130 18570 -1040 18810
rect -800 18570 -710 18810
rect -470 18570 -380 18810
rect -140 18570 -50 18810
rect 190 18570 280 18810
rect 520 18570 610 18810
rect 850 18570 940 18810
rect 1180 18570 1270 18810
rect 1510 18570 1600 18810
rect 1840 18570 1930 18810
rect 2170 18570 2260 18810
rect 2500 18570 2590 18810
rect 2830 18570 2920 18810
rect 3160 18570 3250 18810
rect 3490 18570 3580 18810
rect 3820 18570 3910 18810
rect 4150 18570 4240 18810
rect 4480 18570 4570 18810
rect 4810 18570 4900 18810
rect 5140 18570 5230 18810
rect 5470 18570 5560 18810
rect 5800 18570 5890 18810
rect 6130 18570 6220 18810
rect 6460 18570 6550 18810
rect 6790 18570 6880 18810
rect 7120 18570 7260 18810
rect -4980 18480 7260 18570
rect -4980 18240 -4670 18480
rect -4430 18240 -4340 18480
rect -4100 18240 -4010 18480
rect -3770 18240 -3680 18480
rect -3440 18240 -3350 18480
rect -3110 18240 -3020 18480
rect -2780 18240 -2690 18480
rect -2450 18240 -2360 18480
rect -2120 18240 -2030 18480
rect -1790 18240 -1700 18480
rect -1460 18240 -1370 18480
rect -1130 18240 -1040 18480
rect -800 18240 -710 18480
rect -470 18240 -380 18480
rect -140 18240 -50 18480
rect 190 18240 280 18480
rect 520 18240 610 18480
rect 850 18240 940 18480
rect 1180 18240 1270 18480
rect 1510 18240 1600 18480
rect 1840 18240 1930 18480
rect 2170 18240 2260 18480
rect 2500 18240 2590 18480
rect 2830 18240 2920 18480
rect 3160 18240 3250 18480
rect 3490 18240 3580 18480
rect 3820 18240 3910 18480
rect 4150 18240 4240 18480
rect 4480 18240 4570 18480
rect 4810 18240 4900 18480
rect 5140 18240 5230 18480
rect 5470 18240 5560 18480
rect 5800 18240 5890 18480
rect 6130 18240 6220 18480
rect 6460 18240 6550 18480
rect 6790 18240 6880 18480
rect 7120 18240 7260 18480
rect -4980 18150 7260 18240
rect -4980 17910 -4670 18150
rect -4430 17910 -4340 18150
rect -4100 17910 -4010 18150
rect -3770 17910 -3680 18150
rect -3440 17910 -3350 18150
rect -3110 17910 -3020 18150
rect -2780 17910 -2690 18150
rect -2450 17910 -2360 18150
rect -2120 17910 -2030 18150
rect -1790 17910 -1700 18150
rect -1460 17910 -1370 18150
rect -1130 17910 -1040 18150
rect -800 17910 -710 18150
rect -470 17910 -380 18150
rect -140 17910 -50 18150
rect 190 17910 280 18150
rect 520 17910 610 18150
rect 850 17910 940 18150
rect 1180 17910 1270 18150
rect 1510 17910 1600 18150
rect 1840 17910 1930 18150
rect 2170 17910 2260 18150
rect 2500 17910 2590 18150
rect 2830 17910 2920 18150
rect 3160 17910 3250 18150
rect 3490 17910 3580 18150
rect 3820 17910 3910 18150
rect 4150 17910 4240 18150
rect 4480 17910 4570 18150
rect 4810 17910 4900 18150
rect 5140 17910 5230 18150
rect 5470 17910 5560 18150
rect 5800 17910 5890 18150
rect 6130 17910 6220 18150
rect 6460 17910 6550 18150
rect 6790 17910 6880 18150
rect 7120 17910 7260 18150
rect -4980 17820 7260 17910
rect -4980 17580 -4670 17820
rect -4430 17580 -4340 17820
rect -4100 17580 -4010 17820
rect -3770 17580 -3680 17820
rect -3440 17580 -3350 17820
rect -3110 17580 -3020 17820
rect -2780 17580 -2690 17820
rect -2450 17580 -2360 17820
rect -2120 17580 -2030 17820
rect -1790 17580 -1700 17820
rect -1460 17580 -1370 17820
rect -1130 17580 -1040 17820
rect -800 17580 -710 17820
rect -470 17580 -380 17820
rect -140 17580 -50 17820
rect 190 17580 280 17820
rect 520 17580 610 17820
rect 850 17580 940 17820
rect 1180 17580 1270 17820
rect 1510 17580 1600 17820
rect 1840 17580 1930 17820
rect 2170 17580 2260 17820
rect 2500 17580 2590 17820
rect 2830 17580 2920 17820
rect 3160 17580 3250 17820
rect 3490 17580 3580 17820
rect 3820 17580 3910 17820
rect 4150 17580 4240 17820
rect 4480 17580 4570 17820
rect 4810 17580 4900 17820
rect 5140 17580 5230 17820
rect 5470 17580 5560 17820
rect 5800 17580 5890 17820
rect 6130 17580 6220 17820
rect 6460 17580 6550 17820
rect 6790 17580 6880 17820
rect 7120 17580 7260 17820
rect -4980 17490 7260 17580
rect -4980 17250 -4670 17490
rect -4430 17250 -4340 17490
rect -4100 17250 -4010 17490
rect -3770 17250 -3680 17490
rect -3440 17250 -3350 17490
rect -3110 17250 -3020 17490
rect -2780 17250 -2690 17490
rect -2450 17250 -2360 17490
rect -2120 17250 -2030 17490
rect -1790 17250 -1700 17490
rect -1460 17250 -1370 17490
rect -1130 17250 -1040 17490
rect -800 17250 -710 17490
rect -470 17250 -380 17490
rect -140 17250 -50 17490
rect 190 17250 280 17490
rect 520 17250 610 17490
rect 850 17250 940 17490
rect 1180 17250 1270 17490
rect 1510 17250 1600 17490
rect 1840 17250 1930 17490
rect 2170 17250 2260 17490
rect 2500 17250 2590 17490
rect 2830 17250 2920 17490
rect 3160 17250 3250 17490
rect 3490 17250 3580 17490
rect 3820 17250 3910 17490
rect 4150 17250 4240 17490
rect 4480 17250 4570 17490
rect 4810 17250 4900 17490
rect 5140 17250 5230 17490
rect 5470 17250 5560 17490
rect 5800 17250 5890 17490
rect 6130 17250 6220 17490
rect 6460 17250 6550 17490
rect 6790 17250 6880 17490
rect 7120 17250 7260 17490
rect -4980 17160 7260 17250
rect -4980 16920 -4670 17160
rect -4430 16920 -4340 17160
rect -4100 16920 -4010 17160
rect -3770 16920 -3680 17160
rect -3440 16920 -3350 17160
rect -3110 16920 -3020 17160
rect -2780 16920 -2690 17160
rect -2450 16920 -2360 17160
rect -2120 16920 -2030 17160
rect -1790 16920 -1700 17160
rect -1460 16920 -1370 17160
rect -1130 16920 -1040 17160
rect -800 16920 -710 17160
rect -470 16920 -380 17160
rect -140 16920 -50 17160
rect 190 16920 280 17160
rect 520 16920 610 17160
rect 850 16920 940 17160
rect 1180 16920 1270 17160
rect 1510 16920 1600 17160
rect 1840 16920 1930 17160
rect 2170 16920 2260 17160
rect 2500 16920 2590 17160
rect 2830 16920 2920 17160
rect 3160 16920 3250 17160
rect 3490 16920 3580 17160
rect 3820 16920 3910 17160
rect 4150 16920 4240 17160
rect 4480 16920 4570 17160
rect 4810 16920 4900 17160
rect 5140 16920 5230 17160
rect 5470 16920 5560 17160
rect 5800 16920 5890 17160
rect 6130 16920 6220 17160
rect 6460 16920 6550 17160
rect 6790 16920 6880 17160
rect 7120 16920 7260 17160
rect -4980 16830 7260 16920
rect -4980 16590 -4670 16830
rect -4430 16590 -4340 16830
rect -4100 16590 -4010 16830
rect -3770 16590 -3680 16830
rect -3440 16590 -3350 16830
rect -3110 16590 -3020 16830
rect -2780 16590 -2690 16830
rect -2450 16590 -2360 16830
rect -2120 16590 -2030 16830
rect -1790 16590 -1700 16830
rect -1460 16590 -1370 16830
rect -1130 16590 -1040 16830
rect -800 16590 -710 16830
rect -470 16590 -380 16830
rect -140 16590 -50 16830
rect 190 16590 280 16830
rect 520 16590 610 16830
rect 850 16590 940 16830
rect 1180 16590 1270 16830
rect 1510 16590 1600 16830
rect 1840 16590 1930 16830
rect 2170 16590 2260 16830
rect 2500 16590 2590 16830
rect 2830 16590 2920 16830
rect 3160 16590 3250 16830
rect 3490 16590 3580 16830
rect 3820 16590 3910 16830
rect 4150 16590 4240 16830
rect 4480 16590 4570 16830
rect 4810 16590 4900 16830
rect 5140 16590 5230 16830
rect 5470 16590 5560 16830
rect 5800 16590 5890 16830
rect 6130 16590 6220 16830
rect 6460 16590 6550 16830
rect 6790 16590 6880 16830
rect 7120 16590 7260 16830
rect -4980 16500 7260 16590
rect -4980 16260 -4670 16500
rect -4430 16260 -4340 16500
rect -4100 16260 -4010 16500
rect -3770 16260 -3680 16500
rect -3440 16260 -3350 16500
rect -3110 16260 -3020 16500
rect -2780 16260 -2690 16500
rect -2450 16260 -2360 16500
rect -2120 16260 -2030 16500
rect -1790 16260 -1700 16500
rect -1460 16260 -1370 16500
rect -1130 16260 -1040 16500
rect -800 16260 -710 16500
rect -470 16260 -380 16500
rect -140 16260 -50 16500
rect 190 16260 280 16500
rect 520 16260 610 16500
rect 850 16260 940 16500
rect 1180 16260 1270 16500
rect 1510 16260 1600 16500
rect 1840 16260 1930 16500
rect 2170 16260 2260 16500
rect 2500 16260 2590 16500
rect 2830 16260 2920 16500
rect 3160 16260 3250 16500
rect 3490 16260 3580 16500
rect 3820 16260 3910 16500
rect 4150 16260 4240 16500
rect 4480 16260 4570 16500
rect 4810 16260 4900 16500
rect 5140 16260 5230 16500
rect 5470 16260 5560 16500
rect 5800 16260 5890 16500
rect 6130 16260 6220 16500
rect 6460 16260 6550 16500
rect 6790 16260 6880 16500
rect 7120 16260 7260 16500
rect -4980 16170 7260 16260
rect -4980 15930 -4670 16170
rect -4430 15930 -4340 16170
rect -4100 15930 -4010 16170
rect -3770 15930 -3680 16170
rect -3440 15930 -3350 16170
rect -3110 15930 -3020 16170
rect -2780 15930 -2690 16170
rect -2450 15930 -2360 16170
rect -2120 15930 -2030 16170
rect -1790 15930 -1700 16170
rect -1460 15930 -1370 16170
rect -1130 15930 -1040 16170
rect -800 15930 -710 16170
rect -470 15930 -380 16170
rect -140 15930 -50 16170
rect 190 15930 280 16170
rect 520 15930 610 16170
rect 850 15930 940 16170
rect 1180 15930 1270 16170
rect 1510 15930 1600 16170
rect 1840 15930 1930 16170
rect 2170 15930 2260 16170
rect 2500 15930 2590 16170
rect 2830 15930 2920 16170
rect 3160 15930 3250 16170
rect 3490 15930 3580 16170
rect 3820 15930 3910 16170
rect 4150 15930 4240 16170
rect 4480 15930 4570 16170
rect 4810 15930 4900 16170
rect 5140 15930 5230 16170
rect 5470 15930 5560 16170
rect 5800 15930 5890 16170
rect 6130 15930 6220 16170
rect 6460 15930 6550 16170
rect 6790 15930 6880 16170
rect 7120 15930 7260 16170
rect -4980 15840 7260 15930
rect -4980 15600 -4670 15840
rect -4430 15600 -4340 15840
rect -4100 15600 -4010 15840
rect -3770 15600 -3680 15840
rect -3440 15600 -3350 15840
rect -3110 15600 -3020 15840
rect -2780 15600 -2690 15840
rect -2450 15600 -2360 15840
rect -2120 15600 -2030 15840
rect -1790 15600 -1700 15840
rect -1460 15600 -1370 15840
rect -1130 15600 -1040 15840
rect -800 15600 -710 15840
rect -470 15600 -380 15840
rect -140 15600 -50 15840
rect 190 15600 280 15840
rect 520 15600 610 15840
rect 850 15600 940 15840
rect 1180 15600 1270 15840
rect 1510 15600 1600 15840
rect 1840 15600 1930 15840
rect 2170 15600 2260 15840
rect 2500 15600 2590 15840
rect 2830 15600 2920 15840
rect 3160 15600 3250 15840
rect 3490 15600 3580 15840
rect 3820 15600 3910 15840
rect 4150 15600 4240 15840
rect 4480 15600 4570 15840
rect 4810 15600 4900 15840
rect 5140 15600 5230 15840
rect 5470 15600 5560 15840
rect 5800 15600 5890 15840
rect 6130 15600 6220 15840
rect 6460 15600 6550 15840
rect 6790 15600 6880 15840
rect 7120 15600 7260 15840
rect -4980 15510 7260 15600
rect -4980 15270 -4670 15510
rect -4430 15270 -4340 15510
rect -4100 15270 -4010 15510
rect -3770 15270 -3680 15510
rect -3440 15270 -3350 15510
rect -3110 15270 -3020 15510
rect -2780 15270 -2690 15510
rect -2450 15270 -2360 15510
rect -2120 15270 -2030 15510
rect -1790 15270 -1700 15510
rect -1460 15270 -1370 15510
rect -1130 15270 -1040 15510
rect -800 15270 -710 15510
rect -470 15270 -380 15510
rect -140 15270 -50 15510
rect 190 15270 280 15510
rect 520 15270 610 15510
rect 850 15270 940 15510
rect 1180 15270 1270 15510
rect 1510 15270 1600 15510
rect 1840 15270 1930 15510
rect 2170 15270 2260 15510
rect 2500 15270 2590 15510
rect 2830 15270 2920 15510
rect 3160 15270 3250 15510
rect 3490 15270 3580 15510
rect 3820 15270 3910 15510
rect 4150 15270 4240 15510
rect 4480 15270 4570 15510
rect 4810 15270 4900 15510
rect 5140 15270 5230 15510
rect 5470 15270 5560 15510
rect 5800 15270 5890 15510
rect 6130 15270 6220 15510
rect 6460 15270 6550 15510
rect 6790 15270 6880 15510
rect 7120 15270 7260 15510
rect -4980 15180 7260 15270
rect -4980 14940 -4670 15180
rect -4430 14940 -4340 15180
rect -4100 14940 -4010 15180
rect -3770 14940 -3680 15180
rect -3440 14940 -3350 15180
rect -3110 14940 -3020 15180
rect -2780 14940 -2690 15180
rect -2450 14940 -2360 15180
rect -2120 14940 -2030 15180
rect -1790 14940 -1700 15180
rect -1460 14940 -1370 15180
rect -1130 14940 -1040 15180
rect -800 14940 -710 15180
rect -470 14940 -380 15180
rect -140 14940 -50 15180
rect 190 14940 280 15180
rect 520 14940 610 15180
rect 850 14940 940 15180
rect 1180 14940 1270 15180
rect 1510 14940 1600 15180
rect 1840 14940 1930 15180
rect 2170 14940 2260 15180
rect 2500 14940 2590 15180
rect 2830 14940 2920 15180
rect 3160 14940 3250 15180
rect 3490 14940 3580 15180
rect 3820 14940 3910 15180
rect 4150 14940 4240 15180
rect 4480 14940 4570 15180
rect 4810 14940 4900 15180
rect 5140 14940 5230 15180
rect 5470 14940 5560 15180
rect 5800 14940 5890 15180
rect 6130 14940 6220 15180
rect 6460 14940 6550 15180
rect 6790 14940 6880 15180
rect 7120 14940 7260 15180
rect -4980 14850 7260 14940
rect -4980 14610 -4670 14850
rect -4430 14610 -4340 14850
rect -4100 14610 -4010 14850
rect -3770 14610 -3680 14850
rect -3440 14610 -3350 14850
rect -3110 14610 -3020 14850
rect -2780 14610 -2690 14850
rect -2450 14610 -2360 14850
rect -2120 14610 -2030 14850
rect -1790 14610 -1700 14850
rect -1460 14610 -1370 14850
rect -1130 14610 -1040 14850
rect -800 14610 -710 14850
rect -470 14610 -380 14850
rect -140 14610 -50 14850
rect 190 14610 280 14850
rect 520 14610 610 14850
rect 850 14610 940 14850
rect 1180 14610 1270 14850
rect 1510 14610 1600 14850
rect 1840 14610 1930 14850
rect 2170 14610 2260 14850
rect 2500 14610 2590 14850
rect 2830 14610 2920 14850
rect 3160 14610 3250 14850
rect 3490 14610 3580 14850
rect 3820 14610 3910 14850
rect 4150 14610 4240 14850
rect 4480 14610 4570 14850
rect 4810 14610 4900 14850
rect 5140 14610 5230 14850
rect 5470 14610 5560 14850
rect 5800 14610 5890 14850
rect 6130 14610 6220 14850
rect 6460 14610 6550 14850
rect 6790 14610 6880 14850
rect 7120 14610 7260 14850
rect -4980 14520 7260 14610
rect -4980 14280 -4670 14520
rect -4430 14280 -4340 14520
rect -4100 14280 -4010 14520
rect -3770 14280 -3680 14520
rect -3440 14280 -3350 14520
rect -3110 14280 -3020 14520
rect -2780 14280 -2690 14520
rect -2450 14280 -2360 14520
rect -2120 14280 -2030 14520
rect -1790 14280 -1700 14520
rect -1460 14280 -1370 14520
rect -1130 14280 -1040 14520
rect -800 14280 -710 14520
rect -470 14280 -380 14520
rect -140 14280 -50 14520
rect 190 14280 280 14520
rect 520 14280 610 14520
rect 850 14280 940 14520
rect 1180 14280 1270 14520
rect 1510 14280 1600 14520
rect 1840 14280 1930 14520
rect 2170 14280 2260 14520
rect 2500 14280 2590 14520
rect 2830 14280 2920 14520
rect 3160 14280 3250 14520
rect 3490 14280 3580 14520
rect 3820 14280 3910 14520
rect 4150 14280 4240 14520
rect 4480 14280 4570 14520
rect 4810 14280 4900 14520
rect 5140 14280 5230 14520
rect 5470 14280 5560 14520
rect 5800 14280 5890 14520
rect 6130 14280 6220 14520
rect 6460 14280 6550 14520
rect 6790 14280 6880 14520
rect 7120 14280 7260 14520
rect -4980 14190 7260 14280
rect -4980 13950 -4670 14190
rect -4430 13950 -4340 14190
rect -4100 13950 -4010 14190
rect -3770 13950 -3680 14190
rect -3440 13950 -3350 14190
rect -3110 13950 -3020 14190
rect -2780 13950 -2690 14190
rect -2450 13950 -2360 14190
rect -2120 13950 -2030 14190
rect -1790 13950 -1700 14190
rect -1460 13950 -1370 14190
rect -1130 13950 -1040 14190
rect -800 13950 -710 14190
rect -470 13950 -380 14190
rect -140 13950 -50 14190
rect 190 13950 280 14190
rect 520 13950 610 14190
rect 850 13950 940 14190
rect 1180 13950 1270 14190
rect 1510 13950 1600 14190
rect 1840 13950 1930 14190
rect 2170 13950 2260 14190
rect 2500 13950 2590 14190
rect 2830 13950 2920 14190
rect 3160 13950 3250 14190
rect 3490 13950 3580 14190
rect 3820 13950 3910 14190
rect 4150 13950 4240 14190
rect 4480 13950 4570 14190
rect 4810 13950 4900 14190
rect 5140 13950 5230 14190
rect 5470 13950 5560 14190
rect 5800 13950 5890 14190
rect 6130 13950 6220 14190
rect 6460 13950 6550 14190
rect 6790 13950 6880 14190
rect 7120 13950 7260 14190
rect -4980 13860 7260 13950
rect -4980 13620 -4670 13860
rect -4430 13620 -4340 13860
rect -4100 13620 -4010 13860
rect -3770 13620 -3680 13860
rect -3440 13620 -3350 13860
rect -3110 13620 -3020 13860
rect -2780 13620 -2690 13860
rect -2450 13620 -2360 13860
rect -2120 13620 -2030 13860
rect -1790 13620 -1700 13860
rect -1460 13620 -1370 13860
rect -1130 13620 -1040 13860
rect -800 13620 -710 13860
rect -470 13620 -380 13860
rect -140 13620 -50 13860
rect 190 13620 280 13860
rect 520 13620 610 13860
rect 850 13620 940 13860
rect 1180 13620 1270 13860
rect 1510 13620 1600 13860
rect 1840 13620 1930 13860
rect 2170 13620 2260 13860
rect 2500 13620 2590 13860
rect 2830 13620 2920 13860
rect 3160 13620 3250 13860
rect 3490 13620 3580 13860
rect 3820 13620 3910 13860
rect 4150 13620 4240 13860
rect 4480 13620 4570 13860
rect 4810 13620 4900 13860
rect 5140 13620 5230 13860
rect 5470 13620 5560 13860
rect 5800 13620 5890 13860
rect 6130 13620 6220 13860
rect 6460 13620 6550 13860
rect 6790 13620 6880 13860
rect 7120 13620 7260 13860
rect -4980 13530 7260 13620
rect -4980 13290 -4670 13530
rect -4430 13290 -4340 13530
rect -4100 13290 -4010 13530
rect -3770 13290 -3680 13530
rect -3440 13290 -3350 13530
rect -3110 13290 -3020 13530
rect -2780 13290 -2690 13530
rect -2450 13290 -2360 13530
rect -2120 13290 -2030 13530
rect -1790 13290 -1700 13530
rect -1460 13290 -1370 13530
rect -1130 13290 -1040 13530
rect -800 13290 -710 13530
rect -470 13290 -380 13530
rect -140 13290 -50 13530
rect 190 13290 280 13530
rect 520 13290 610 13530
rect 850 13290 940 13530
rect 1180 13290 1270 13530
rect 1510 13290 1600 13530
rect 1840 13290 1930 13530
rect 2170 13290 2260 13530
rect 2500 13290 2590 13530
rect 2830 13290 2920 13530
rect 3160 13290 3250 13530
rect 3490 13290 3580 13530
rect 3820 13290 3910 13530
rect 4150 13290 4240 13530
rect 4480 13290 4570 13530
rect 4810 13290 4900 13530
rect 5140 13290 5230 13530
rect 5470 13290 5560 13530
rect 5800 13290 5890 13530
rect 6130 13290 6220 13530
rect 6460 13290 6550 13530
rect 6790 13290 6880 13530
rect 7120 13290 7260 13530
rect -4980 13200 7260 13290
rect -4980 12960 -4670 13200
rect -4430 12960 -4340 13200
rect -4100 12960 -4010 13200
rect -3770 12960 -3680 13200
rect -3440 12960 -3350 13200
rect -3110 12960 -3020 13200
rect -2780 12960 -2690 13200
rect -2450 12960 -2360 13200
rect -2120 12960 -2030 13200
rect -1790 12960 -1700 13200
rect -1460 12960 -1370 13200
rect -1130 12960 -1040 13200
rect -800 12960 -710 13200
rect -470 12960 -380 13200
rect -140 12960 -50 13200
rect 190 12960 280 13200
rect 520 12960 610 13200
rect 850 12960 940 13200
rect 1180 12960 1270 13200
rect 1510 12960 1600 13200
rect 1840 12960 1930 13200
rect 2170 12960 2260 13200
rect 2500 12960 2590 13200
rect 2830 12960 2920 13200
rect 3160 12960 3250 13200
rect 3490 12960 3580 13200
rect 3820 12960 3910 13200
rect 4150 12960 4240 13200
rect 4480 12960 4570 13200
rect 4810 12960 4900 13200
rect 5140 12960 5230 13200
rect 5470 12960 5560 13200
rect 5800 12960 5890 13200
rect 6130 12960 6220 13200
rect 6460 12960 6550 13200
rect 6790 12960 6880 13200
rect 7120 12960 7260 13200
rect -4980 12870 7260 12960
rect -4980 12630 -4670 12870
rect -4430 12630 -4340 12870
rect -4100 12630 -4010 12870
rect -3770 12630 -3680 12870
rect -3440 12630 -3350 12870
rect -3110 12630 -3020 12870
rect -2780 12630 -2690 12870
rect -2450 12630 -2360 12870
rect -2120 12630 -2030 12870
rect -1790 12630 -1700 12870
rect -1460 12630 -1370 12870
rect -1130 12630 -1040 12870
rect -800 12630 -710 12870
rect -470 12630 -380 12870
rect -140 12630 -50 12870
rect 190 12630 280 12870
rect 520 12630 610 12870
rect 850 12630 940 12870
rect 1180 12630 1270 12870
rect 1510 12630 1600 12870
rect 1840 12630 1930 12870
rect 2170 12630 2260 12870
rect 2500 12630 2590 12870
rect 2830 12630 2920 12870
rect 3160 12630 3250 12870
rect 3490 12630 3580 12870
rect 3820 12630 3910 12870
rect 4150 12630 4240 12870
rect 4480 12630 4570 12870
rect 4810 12630 4900 12870
rect 5140 12630 5230 12870
rect 5470 12630 5560 12870
rect 5800 12630 5890 12870
rect 6130 12630 6220 12870
rect 6460 12630 6550 12870
rect 6790 12630 6880 12870
rect 7120 12630 7260 12870
rect -4980 12540 7260 12630
rect -4980 12300 -4670 12540
rect -4430 12300 -4340 12540
rect -4100 12300 -4010 12540
rect -3770 12300 -3680 12540
rect -3440 12300 -3350 12540
rect -3110 12300 -3020 12540
rect -2780 12300 -2690 12540
rect -2450 12300 -2360 12540
rect -2120 12300 -2030 12540
rect -1790 12300 -1700 12540
rect -1460 12300 -1370 12540
rect -1130 12300 -1040 12540
rect -800 12300 -710 12540
rect -470 12300 -380 12540
rect -140 12300 -50 12540
rect 190 12300 280 12540
rect 520 12300 610 12540
rect 850 12300 940 12540
rect 1180 12300 1270 12540
rect 1510 12300 1600 12540
rect 1840 12300 1930 12540
rect 2170 12300 2260 12540
rect 2500 12300 2590 12540
rect 2830 12300 2920 12540
rect 3160 12300 3250 12540
rect 3490 12300 3580 12540
rect 3820 12300 3910 12540
rect 4150 12300 4240 12540
rect 4480 12300 4570 12540
rect 4810 12300 4900 12540
rect 5140 12300 5230 12540
rect 5470 12300 5560 12540
rect 5800 12300 5890 12540
rect 6130 12300 6220 12540
rect 6460 12300 6550 12540
rect 6790 12300 6880 12540
rect 7120 12300 7260 12540
rect -4980 12210 7260 12300
rect -4980 11970 -4670 12210
rect -4430 11970 -4340 12210
rect -4100 11970 -4010 12210
rect -3770 11970 -3680 12210
rect -3440 11970 -3350 12210
rect -3110 11970 -3020 12210
rect -2780 11970 -2690 12210
rect -2450 11970 -2360 12210
rect -2120 11970 -2030 12210
rect -1790 11970 -1700 12210
rect -1460 11970 -1370 12210
rect -1130 11970 -1040 12210
rect -800 11970 -710 12210
rect -470 11970 -380 12210
rect -140 11970 -50 12210
rect 190 11970 280 12210
rect 520 11970 610 12210
rect 850 11970 940 12210
rect 1180 11970 1270 12210
rect 1510 11970 1600 12210
rect 1840 11970 1930 12210
rect 2170 11970 2260 12210
rect 2500 11970 2590 12210
rect 2830 11970 2920 12210
rect 3160 11970 3250 12210
rect 3490 11970 3580 12210
rect 3820 11970 3910 12210
rect 4150 11970 4240 12210
rect 4480 11970 4570 12210
rect 4810 11970 4900 12210
rect 5140 11970 5230 12210
rect 5470 11970 5560 12210
rect 5800 11970 5890 12210
rect 6130 11970 6220 12210
rect 6460 11970 6550 12210
rect 6790 11970 6880 12210
rect 7120 11970 7260 12210
rect -4980 11880 7260 11970
rect -4980 11640 -4670 11880
rect -4430 11640 -4340 11880
rect -4100 11640 -4010 11880
rect -3770 11640 -3680 11880
rect -3440 11640 -3350 11880
rect -3110 11640 -3020 11880
rect -2780 11640 -2690 11880
rect -2450 11640 -2360 11880
rect -2120 11640 -2030 11880
rect -1790 11640 -1700 11880
rect -1460 11640 -1370 11880
rect -1130 11640 -1040 11880
rect -800 11640 -710 11880
rect -470 11640 -380 11880
rect -140 11640 -50 11880
rect 190 11640 280 11880
rect 520 11640 610 11880
rect 850 11640 940 11880
rect 1180 11640 1270 11880
rect 1510 11640 1600 11880
rect 1840 11640 1930 11880
rect 2170 11640 2260 11880
rect 2500 11640 2590 11880
rect 2830 11640 2920 11880
rect 3160 11640 3250 11880
rect 3490 11640 3580 11880
rect 3820 11640 3910 11880
rect 4150 11640 4240 11880
rect 4480 11640 4570 11880
rect 4810 11640 4900 11880
rect 5140 11640 5230 11880
rect 5470 11640 5560 11880
rect 5800 11640 5890 11880
rect 6130 11640 6220 11880
rect 6460 11640 6550 11880
rect 6790 11640 6880 11880
rect 7120 11640 7260 11880
rect -4980 11550 7260 11640
rect -4980 11310 -4670 11550
rect -4430 11310 -4340 11550
rect -4100 11310 -4010 11550
rect -3770 11310 -3680 11550
rect -3440 11310 -3350 11550
rect -3110 11310 -3020 11550
rect -2780 11310 -2690 11550
rect -2450 11310 -2360 11550
rect -2120 11310 -2030 11550
rect -1790 11310 -1700 11550
rect -1460 11310 -1370 11550
rect -1130 11310 -1040 11550
rect -800 11310 -710 11550
rect -470 11310 -380 11550
rect -140 11310 -50 11550
rect 190 11310 280 11550
rect 520 11310 610 11550
rect 850 11310 940 11550
rect 1180 11310 1270 11550
rect 1510 11310 1600 11550
rect 1840 11310 1930 11550
rect 2170 11310 2260 11550
rect 2500 11310 2590 11550
rect 2830 11310 2920 11550
rect 3160 11310 3250 11550
rect 3490 11310 3580 11550
rect 3820 11310 3910 11550
rect 4150 11310 4240 11550
rect 4480 11310 4570 11550
rect 4810 11310 4900 11550
rect 5140 11310 5230 11550
rect 5470 11310 5560 11550
rect 5800 11310 5890 11550
rect 6130 11310 6220 11550
rect 6460 11310 6550 11550
rect 6790 11310 6880 11550
rect 7120 11310 7260 11550
rect -4980 11220 7260 11310
rect -4980 10980 -4670 11220
rect -4430 10980 -4340 11220
rect -4100 10980 -4010 11220
rect -3770 10980 -3680 11220
rect -3440 10980 -3350 11220
rect -3110 10980 -3020 11220
rect -2780 10980 -2690 11220
rect -2450 10980 -2360 11220
rect -2120 10980 -2030 11220
rect -1790 10980 -1700 11220
rect -1460 10980 -1370 11220
rect -1130 10980 -1040 11220
rect -800 10980 -710 11220
rect -470 10980 -380 11220
rect -140 10980 -50 11220
rect 190 10980 280 11220
rect 520 10980 610 11220
rect 850 10980 940 11220
rect 1180 10980 1270 11220
rect 1510 10980 1600 11220
rect 1840 10980 1930 11220
rect 2170 10980 2260 11220
rect 2500 10980 2590 11220
rect 2830 10980 2920 11220
rect 3160 10980 3250 11220
rect 3490 10980 3580 11220
rect 3820 10980 3910 11220
rect 4150 10980 4240 11220
rect 4480 10980 4570 11220
rect 4810 10980 4900 11220
rect 5140 10980 5230 11220
rect 5470 10980 5560 11220
rect 5800 10980 5890 11220
rect 6130 10980 6220 11220
rect 6460 10980 6550 11220
rect 6790 10980 6880 11220
rect 7120 10980 7260 11220
rect -4980 10890 7260 10980
rect -4980 10650 -4670 10890
rect -4430 10650 -4340 10890
rect -4100 10650 -4010 10890
rect -3770 10650 -3680 10890
rect -3440 10650 -3350 10890
rect -3110 10650 -3020 10890
rect -2780 10650 -2690 10890
rect -2450 10650 -2360 10890
rect -2120 10650 -2030 10890
rect -1790 10650 -1700 10890
rect -1460 10650 -1370 10890
rect -1130 10650 -1040 10890
rect -800 10650 -710 10890
rect -470 10650 -380 10890
rect -140 10650 -50 10890
rect 190 10650 280 10890
rect 520 10650 610 10890
rect 850 10650 940 10890
rect 1180 10650 1270 10890
rect 1510 10650 1600 10890
rect 1840 10650 1930 10890
rect 2170 10650 2260 10890
rect 2500 10650 2590 10890
rect 2830 10650 2920 10890
rect 3160 10650 3250 10890
rect 3490 10650 3580 10890
rect 3820 10650 3910 10890
rect 4150 10650 4240 10890
rect 4480 10650 4570 10890
rect 4810 10650 4900 10890
rect 5140 10650 5230 10890
rect 5470 10650 5560 10890
rect 5800 10650 5890 10890
rect 6130 10650 6220 10890
rect 6460 10650 6550 10890
rect 6790 10650 6880 10890
rect 7120 10650 7260 10890
rect -4980 10560 7260 10650
rect -4980 10320 -4670 10560
rect -4430 10320 -4340 10560
rect -4100 10320 -4010 10560
rect -3770 10320 -3680 10560
rect -3440 10320 -3350 10560
rect -3110 10320 -3020 10560
rect -2780 10320 -2690 10560
rect -2450 10320 -2360 10560
rect -2120 10320 -2030 10560
rect -1790 10320 -1700 10560
rect -1460 10320 -1370 10560
rect -1130 10320 -1040 10560
rect -800 10320 -710 10560
rect -470 10320 -380 10560
rect -140 10320 -50 10560
rect 190 10320 280 10560
rect 520 10320 610 10560
rect 850 10320 940 10560
rect 1180 10320 1270 10560
rect 1510 10320 1600 10560
rect 1840 10320 1930 10560
rect 2170 10320 2260 10560
rect 2500 10320 2590 10560
rect 2830 10320 2920 10560
rect 3160 10320 3250 10560
rect 3490 10320 3580 10560
rect 3820 10320 3910 10560
rect 4150 10320 4240 10560
rect 4480 10320 4570 10560
rect 4810 10320 4900 10560
rect 5140 10320 5230 10560
rect 5470 10320 5560 10560
rect 5800 10320 5890 10560
rect 6130 10320 6220 10560
rect 6460 10320 6550 10560
rect 6790 10320 6880 10560
rect 7120 10320 7260 10560
rect -4980 10230 7260 10320
rect -4980 9990 -4670 10230
rect -4430 9990 -4340 10230
rect -4100 9990 -4010 10230
rect -3770 9990 -3680 10230
rect -3440 9990 -3350 10230
rect -3110 9990 -3020 10230
rect -2780 9990 -2690 10230
rect -2450 9990 -2360 10230
rect -2120 9990 -2030 10230
rect -1790 9990 -1700 10230
rect -1460 9990 -1370 10230
rect -1130 9990 -1040 10230
rect -800 9990 -710 10230
rect -470 9990 -380 10230
rect -140 9990 -50 10230
rect 190 9990 280 10230
rect 520 9990 610 10230
rect 850 9990 940 10230
rect 1180 9990 1270 10230
rect 1510 9990 1600 10230
rect 1840 9990 1930 10230
rect 2170 9990 2260 10230
rect 2500 9990 2590 10230
rect 2830 9990 2920 10230
rect 3160 9990 3250 10230
rect 3490 9990 3580 10230
rect 3820 9990 3910 10230
rect 4150 9990 4240 10230
rect 4480 9990 4570 10230
rect 4810 9990 4900 10230
rect 5140 9990 5230 10230
rect 5470 9990 5560 10230
rect 5800 9990 5890 10230
rect 6130 9990 6220 10230
rect 6460 9990 6550 10230
rect 6790 9990 6880 10230
rect 7120 9990 7260 10230
rect -4980 9900 7260 9990
rect -4980 9660 -4670 9900
rect -4430 9660 -4340 9900
rect -4100 9660 -4010 9900
rect -3770 9660 -3680 9900
rect -3440 9660 -3350 9900
rect -3110 9660 -3020 9900
rect -2780 9660 -2690 9900
rect -2450 9660 -2360 9900
rect -2120 9660 -2030 9900
rect -1790 9660 -1700 9900
rect -1460 9660 -1370 9900
rect -1130 9660 -1040 9900
rect -800 9660 -710 9900
rect -470 9660 -380 9900
rect -140 9660 -50 9900
rect 190 9660 280 9900
rect 520 9660 610 9900
rect 850 9660 940 9900
rect 1180 9660 1270 9900
rect 1510 9660 1600 9900
rect 1840 9660 1930 9900
rect 2170 9660 2260 9900
rect 2500 9660 2590 9900
rect 2830 9660 2920 9900
rect 3160 9660 3250 9900
rect 3490 9660 3580 9900
rect 3820 9660 3910 9900
rect 4150 9660 4240 9900
rect 4480 9660 4570 9900
rect 4810 9660 4900 9900
rect 5140 9660 5230 9900
rect 5470 9660 5560 9900
rect 5800 9660 5890 9900
rect 6130 9660 6220 9900
rect 6460 9660 6550 9900
rect 6790 9660 6880 9900
rect 7120 9660 7260 9900
rect -4980 9570 7260 9660
rect -4980 9330 -4670 9570
rect -4430 9330 -4340 9570
rect -4100 9330 -4010 9570
rect -3770 9330 -3680 9570
rect -3440 9330 -3350 9570
rect -3110 9330 -3020 9570
rect -2780 9330 -2690 9570
rect -2450 9330 -2360 9570
rect -2120 9330 -2030 9570
rect -1790 9330 -1700 9570
rect -1460 9330 -1370 9570
rect -1130 9330 -1040 9570
rect -800 9330 -710 9570
rect -470 9330 -380 9570
rect -140 9330 -50 9570
rect 190 9330 280 9570
rect 520 9330 610 9570
rect 850 9330 940 9570
rect 1180 9330 1270 9570
rect 1510 9330 1600 9570
rect 1840 9330 1930 9570
rect 2170 9330 2260 9570
rect 2500 9330 2590 9570
rect 2830 9330 2920 9570
rect 3160 9330 3250 9570
rect 3490 9330 3580 9570
rect 3820 9330 3910 9570
rect 4150 9330 4240 9570
rect 4480 9330 4570 9570
rect 4810 9330 4900 9570
rect 5140 9330 5230 9570
rect 5470 9330 5560 9570
rect 5800 9330 5890 9570
rect 6130 9330 6220 9570
rect 6460 9330 6550 9570
rect 6790 9330 6880 9570
rect 7120 9330 7260 9570
rect -4980 9240 7260 9330
rect -4980 9000 -4670 9240
rect -4430 9000 -4340 9240
rect -4100 9000 -4010 9240
rect -3770 9000 -3680 9240
rect -3440 9000 -3350 9240
rect -3110 9000 -3020 9240
rect -2780 9000 -2690 9240
rect -2450 9000 -2360 9240
rect -2120 9000 -2030 9240
rect -1790 9000 -1700 9240
rect -1460 9000 -1370 9240
rect -1130 9000 -1040 9240
rect -800 9000 -710 9240
rect -470 9000 -380 9240
rect -140 9000 -50 9240
rect 190 9000 280 9240
rect 520 9000 610 9240
rect 850 9000 940 9240
rect 1180 9000 1270 9240
rect 1510 9000 1600 9240
rect 1840 9000 1930 9240
rect 2170 9000 2260 9240
rect 2500 9000 2590 9240
rect 2830 9000 2920 9240
rect 3160 9000 3250 9240
rect 3490 9000 3580 9240
rect 3820 9000 3910 9240
rect 4150 9000 4240 9240
rect 4480 9000 4570 9240
rect 4810 9000 4900 9240
rect 5140 9000 5230 9240
rect 5470 9000 5560 9240
rect 5800 9000 5890 9240
rect 6130 9000 6220 9240
rect 6460 9000 6550 9240
rect 6790 9000 6880 9240
rect 7120 9000 7260 9240
rect -4980 8870 7260 9000
rect 7640 20790 19880 21110
rect 7640 20550 7780 20790
rect 8020 20550 8110 20790
rect 8350 20550 8440 20790
rect 8680 20550 8770 20790
rect 9010 20550 9100 20790
rect 9340 20550 9430 20790
rect 9670 20550 9760 20790
rect 10000 20550 10090 20790
rect 10330 20550 10420 20790
rect 10660 20550 10750 20790
rect 10990 20550 11080 20790
rect 11320 20550 11410 20790
rect 11650 20550 11740 20790
rect 11980 20550 12070 20790
rect 12310 20550 12400 20790
rect 12640 20550 12730 20790
rect 12970 20550 13060 20790
rect 13300 20550 13390 20790
rect 13630 20550 13720 20790
rect 13960 20550 14050 20790
rect 14290 20550 14380 20790
rect 14620 20550 14710 20790
rect 14950 20550 15040 20790
rect 15280 20550 15370 20790
rect 15610 20550 15700 20790
rect 15940 20550 16030 20790
rect 16270 20550 16360 20790
rect 16600 20550 16690 20790
rect 16930 20550 17020 20790
rect 17260 20550 17350 20790
rect 17590 20550 17680 20790
rect 17920 20550 18010 20790
rect 18250 20550 18340 20790
rect 18580 20550 18670 20790
rect 18910 20550 19000 20790
rect 19240 20550 19330 20790
rect 19570 20550 19880 20790
rect 7640 20460 19880 20550
rect 7640 20220 7780 20460
rect 8020 20220 8110 20460
rect 8350 20220 8440 20460
rect 8680 20220 8770 20460
rect 9010 20220 9100 20460
rect 9340 20220 9430 20460
rect 9670 20220 9760 20460
rect 10000 20220 10090 20460
rect 10330 20220 10420 20460
rect 10660 20220 10750 20460
rect 10990 20220 11080 20460
rect 11320 20220 11410 20460
rect 11650 20220 11740 20460
rect 11980 20220 12070 20460
rect 12310 20220 12400 20460
rect 12640 20220 12730 20460
rect 12970 20220 13060 20460
rect 13300 20220 13390 20460
rect 13630 20220 13720 20460
rect 13960 20220 14050 20460
rect 14290 20220 14380 20460
rect 14620 20220 14710 20460
rect 14950 20220 15040 20460
rect 15280 20220 15370 20460
rect 15610 20220 15700 20460
rect 15940 20220 16030 20460
rect 16270 20220 16360 20460
rect 16600 20220 16690 20460
rect 16930 20220 17020 20460
rect 17260 20220 17350 20460
rect 17590 20220 17680 20460
rect 17920 20220 18010 20460
rect 18250 20220 18340 20460
rect 18580 20220 18670 20460
rect 18910 20220 19000 20460
rect 19240 20220 19330 20460
rect 19570 20220 19880 20460
rect 7640 20130 19880 20220
rect 7640 19890 7780 20130
rect 8020 19890 8110 20130
rect 8350 19890 8440 20130
rect 8680 19890 8770 20130
rect 9010 19890 9100 20130
rect 9340 19890 9430 20130
rect 9670 19890 9760 20130
rect 10000 19890 10090 20130
rect 10330 19890 10420 20130
rect 10660 19890 10750 20130
rect 10990 19890 11080 20130
rect 11320 19890 11410 20130
rect 11650 19890 11740 20130
rect 11980 19890 12070 20130
rect 12310 19890 12400 20130
rect 12640 19890 12730 20130
rect 12970 19890 13060 20130
rect 13300 19890 13390 20130
rect 13630 19890 13720 20130
rect 13960 19890 14050 20130
rect 14290 19890 14380 20130
rect 14620 19890 14710 20130
rect 14950 19890 15040 20130
rect 15280 19890 15370 20130
rect 15610 19890 15700 20130
rect 15940 19890 16030 20130
rect 16270 19890 16360 20130
rect 16600 19890 16690 20130
rect 16930 19890 17020 20130
rect 17260 19890 17350 20130
rect 17590 19890 17680 20130
rect 17920 19890 18010 20130
rect 18250 19890 18340 20130
rect 18580 19890 18670 20130
rect 18910 19890 19000 20130
rect 19240 19890 19330 20130
rect 19570 19890 19880 20130
rect 7640 19800 19880 19890
rect 7640 19560 7780 19800
rect 8020 19560 8110 19800
rect 8350 19560 8440 19800
rect 8680 19560 8770 19800
rect 9010 19560 9100 19800
rect 9340 19560 9430 19800
rect 9670 19560 9760 19800
rect 10000 19560 10090 19800
rect 10330 19560 10420 19800
rect 10660 19560 10750 19800
rect 10990 19560 11080 19800
rect 11320 19560 11410 19800
rect 11650 19560 11740 19800
rect 11980 19560 12070 19800
rect 12310 19560 12400 19800
rect 12640 19560 12730 19800
rect 12970 19560 13060 19800
rect 13300 19560 13390 19800
rect 13630 19560 13720 19800
rect 13960 19560 14050 19800
rect 14290 19560 14380 19800
rect 14620 19560 14710 19800
rect 14950 19560 15040 19800
rect 15280 19560 15370 19800
rect 15610 19560 15700 19800
rect 15940 19560 16030 19800
rect 16270 19560 16360 19800
rect 16600 19560 16690 19800
rect 16930 19560 17020 19800
rect 17260 19560 17350 19800
rect 17590 19560 17680 19800
rect 17920 19560 18010 19800
rect 18250 19560 18340 19800
rect 18580 19560 18670 19800
rect 18910 19560 19000 19800
rect 19240 19560 19330 19800
rect 19570 19560 19880 19800
rect 7640 19470 19880 19560
rect 7640 19230 7780 19470
rect 8020 19230 8110 19470
rect 8350 19230 8440 19470
rect 8680 19230 8770 19470
rect 9010 19230 9100 19470
rect 9340 19230 9430 19470
rect 9670 19230 9760 19470
rect 10000 19230 10090 19470
rect 10330 19230 10420 19470
rect 10660 19230 10750 19470
rect 10990 19230 11080 19470
rect 11320 19230 11410 19470
rect 11650 19230 11740 19470
rect 11980 19230 12070 19470
rect 12310 19230 12400 19470
rect 12640 19230 12730 19470
rect 12970 19230 13060 19470
rect 13300 19230 13390 19470
rect 13630 19230 13720 19470
rect 13960 19230 14050 19470
rect 14290 19230 14380 19470
rect 14620 19230 14710 19470
rect 14950 19230 15040 19470
rect 15280 19230 15370 19470
rect 15610 19230 15700 19470
rect 15940 19230 16030 19470
rect 16270 19230 16360 19470
rect 16600 19230 16690 19470
rect 16930 19230 17020 19470
rect 17260 19230 17350 19470
rect 17590 19230 17680 19470
rect 17920 19230 18010 19470
rect 18250 19230 18340 19470
rect 18580 19230 18670 19470
rect 18910 19230 19000 19470
rect 19240 19230 19330 19470
rect 19570 19230 19880 19470
rect 7640 19140 19880 19230
rect 7640 18900 7780 19140
rect 8020 18900 8110 19140
rect 8350 18900 8440 19140
rect 8680 18900 8770 19140
rect 9010 18900 9100 19140
rect 9340 18900 9430 19140
rect 9670 18900 9760 19140
rect 10000 18900 10090 19140
rect 10330 18900 10420 19140
rect 10660 18900 10750 19140
rect 10990 18900 11080 19140
rect 11320 18900 11410 19140
rect 11650 18900 11740 19140
rect 11980 18900 12070 19140
rect 12310 18900 12400 19140
rect 12640 18900 12730 19140
rect 12970 18900 13060 19140
rect 13300 18900 13390 19140
rect 13630 18900 13720 19140
rect 13960 18900 14050 19140
rect 14290 18900 14380 19140
rect 14620 18900 14710 19140
rect 14950 18900 15040 19140
rect 15280 18900 15370 19140
rect 15610 18900 15700 19140
rect 15940 18900 16030 19140
rect 16270 18900 16360 19140
rect 16600 18900 16690 19140
rect 16930 18900 17020 19140
rect 17260 18900 17350 19140
rect 17590 18900 17680 19140
rect 17920 18900 18010 19140
rect 18250 18900 18340 19140
rect 18580 18900 18670 19140
rect 18910 18900 19000 19140
rect 19240 18900 19330 19140
rect 19570 18900 19880 19140
rect 7640 18810 19880 18900
rect 7640 18570 7780 18810
rect 8020 18570 8110 18810
rect 8350 18570 8440 18810
rect 8680 18570 8770 18810
rect 9010 18570 9100 18810
rect 9340 18570 9430 18810
rect 9670 18570 9760 18810
rect 10000 18570 10090 18810
rect 10330 18570 10420 18810
rect 10660 18570 10750 18810
rect 10990 18570 11080 18810
rect 11320 18570 11410 18810
rect 11650 18570 11740 18810
rect 11980 18570 12070 18810
rect 12310 18570 12400 18810
rect 12640 18570 12730 18810
rect 12970 18570 13060 18810
rect 13300 18570 13390 18810
rect 13630 18570 13720 18810
rect 13960 18570 14050 18810
rect 14290 18570 14380 18810
rect 14620 18570 14710 18810
rect 14950 18570 15040 18810
rect 15280 18570 15370 18810
rect 15610 18570 15700 18810
rect 15940 18570 16030 18810
rect 16270 18570 16360 18810
rect 16600 18570 16690 18810
rect 16930 18570 17020 18810
rect 17260 18570 17350 18810
rect 17590 18570 17680 18810
rect 17920 18570 18010 18810
rect 18250 18570 18340 18810
rect 18580 18570 18670 18810
rect 18910 18570 19000 18810
rect 19240 18570 19330 18810
rect 19570 18570 19880 18810
rect 7640 18480 19880 18570
rect 7640 18240 7780 18480
rect 8020 18240 8110 18480
rect 8350 18240 8440 18480
rect 8680 18240 8770 18480
rect 9010 18240 9100 18480
rect 9340 18240 9430 18480
rect 9670 18240 9760 18480
rect 10000 18240 10090 18480
rect 10330 18240 10420 18480
rect 10660 18240 10750 18480
rect 10990 18240 11080 18480
rect 11320 18240 11410 18480
rect 11650 18240 11740 18480
rect 11980 18240 12070 18480
rect 12310 18240 12400 18480
rect 12640 18240 12730 18480
rect 12970 18240 13060 18480
rect 13300 18240 13390 18480
rect 13630 18240 13720 18480
rect 13960 18240 14050 18480
rect 14290 18240 14380 18480
rect 14620 18240 14710 18480
rect 14950 18240 15040 18480
rect 15280 18240 15370 18480
rect 15610 18240 15700 18480
rect 15940 18240 16030 18480
rect 16270 18240 16360 18480
rect 16600 18240 16690 18480
rect 16930 18240 17020 18480
rect 17260 18240 17350 18480
rect 17590 18240 17680 18480
rect 17920 18240 18010 18480
rect 18250 18240 18340 18480
rect 18580 18240 18670 18480
rect 18910 18240 19000 18480
rect 19240 18240 19330 18480
rect 19570 18240 19880 18480
rect 7640 18150 19880 18240
rect 7640 17910 7780 18150
rect 8020 17910 8110 18150
rect 8350 17910 8440 18150
rect 8680 17910 8770 18150
rect 9010 17910 9100 18150
rect 9340 17910 9430 18150
rect 9670 17910 9760 18150
rect 10000 17910 10090 18150
rect 10330 17910 10420 18150
rect 10660 17910 10750 18150
rect 10990 17910 11080 18150
rect 11320 17910 11410 18150
rect 11650 17910 11740 18150
rect 11980 17910 12070 18150
rect 12310 17910 12400 18150
rect 12640 17910 12730 18150
rect 12970 17910 13060 18150
rect 13300 17910 13390 18150
rect 13630 17910 13720 18150
rect 13960 17910 14050 18150
rect 14290 17910 14380 18150
rect 14620 17910 14710 18150
rect 14950 17910 15040 18150
rect 15280 17910 15370 18150
rect 15610 17910 15700 18150
rect 15940 17910 16030 18150
rect 16270 17910 16360 18150
rect 16600 17910 16690 18150
rect 16930 17910 17020 18150
rect 17260 17910 17350 18150
rect 17590 17910 17680 18150
rect 17920 17910 18010 18150
rect 18250 17910 18340 18150
rect 18580 17910 18670 18150
rect 18910 17910 19000 18150
rect 19240 17910 19330 18150
rect 19570 17910 19880 18150
rect 7640 17820 19880 17910
rect 7640 17580 7780 17820
rect 8020 17580 8110 17820
rect 8350 17580 8440 17820
rect 8680 17580 8770 17820
rect 9010 17580 9100 17820
rect 9340 17580 9430 17820
rect 9670 17580 9760 17820
rect 10000 17580 10090 17820
rect 10330 17580 10420 17820
rect 10660 17580 10750 17820
rect 10990 17580 11080 17820
rect 11320 17580 11410 17820
rect 11650 17580 11740 17820
rect 11980 17580 12070 17820
rect 12310 17580 12400 17820
rect 12640 17580 12730 17820
rect 12970 17580 13060 17820
rect 13300 17580 13390 17820
rect 13630 17580 13720 17820
rect 13960 17580 14050 17820
rect 14290 17580 14380 17820
rect 14620 17580 14710 17820
rect 14950 17580 15040 17820
rect 15280 17580 15370 17820
rect 15610 17580 15700 17820
rect 15940 17580 16030 17820
rect 16270 17580 16360 17820
rect 16600 17580 16690 17820
rect 16930 17580 17020 17820
rect 17260 17580 17350 17820
rect 17590 17580 17680 17820
rect 17920 17580 18010 17820
rect 18250 17580 18340 17820
rect 18580 17580 18670 17820
rect 18910 17580 19000 17820
rect 19240 17580 19330 17820
rect 19570 17580 19880 17820
rect 7640 17490 19880 17580
rect 7640 17250 7780 17490
rect 8020 17250 8110 17490
rect 8350 17250 8440 17490
rect 8680 17250 8770 17490
rect 9010 17250 9100 17490
rect 9340 17250 9430 17490
rect 9670 17250 9760 17490
rect 10000 17250 10090 17490
rect 10330 17250 10420 17490
rect 10660 17250 10750 17490
rect 10990 17250 11080 17490
rect 11320 17250 11410 17490
rect 11650 17250 11740 17490
rect 11980 17250 12070 17490
rect 12310 17250 12400 17490
rect 12640 17250 12730 17490
rect 12970 17250 13060 17490
rect 13300 17250 13390 17490
rect 13630 17250 13720 17490
rect 13960 17250 14050 17490
rect 14290 17250 14380 17490
rect 14620 17250 14710 17490
rect 14950 17250 15040 17490
rect 15280 17250 15370 17490
rect 15610 17250 15700 17490
rect 15940 17250 16030 17490
rect 16270 17250 16360 17490
rect 16600 17250 16690 17490
rect 16930 17250 17020 17490
rect 17260 17250 17350 17490
rect 17590 17250 17680 17490
rect 17920 17250 18010 17490
rect 18250 17250 18340 17490
rect 18580 17250 18670 17490
rect 18910 17250 19000 17490
rect 19240 17250 19330 17490
rect 19570 17250 19880 17490
rect 7640 17160 19880 17250
rect 7640 16920 7780 17160
rect 8020 16920 8110 17160
rect 8350 16920 8440 17160
rect 8680 16920 8770 17160
rect 9010 16920 9100 17160
rect 9340 16920 9430 17160
rect 9670 16920 9760 17160
rect 10000 16920 10090 17160
rect 10330 16920 10420 17160
rect 10660 16920 10750 17160
rect 10990 16920 11080 17160
rect 11320 16920 11410 17160
rect 11650 16920 11740 17160
rect 11980 16920 12070 17160
rect 12310 16920 12400 17160
rect 12640 16920 12730 17160
rect 12970 16920 13060 17160
rect 13300 16920 13390 17160
rect 13630 16920 13720 17160
rect 13960 16920 14050 17160
rect 14290 16920 14380 17160
rect 14620 16920 14710 17160
rect 14950 16920 15040 17160
rect 15280 16920 15370 17160
rect 15610 16920 15700 17160
rect 15940 16920 16030 17160
rect 16270 16920 16360 17160
rect 16600 16920 16690 17160
rect 16930 16920 17020 17160
rect 17260 16920 17350 17160
rect 17590 16920 17680 17160
rect 17920 16920 18010 17160
rect 18250 16920 18340 17160
rect 18580 16920 18670 17160
rect 18910 16920 19000 17160
rect 19240 16920 19330 17160
rect 19570 16920 19880 17160
rect 7640 16830 19880 16920
rect 7640 16590 7780 16830
rect 8020 16590 8110 16830
rect 8350 16590 8440 16830
rect 8680 16590 8770 16830
rect 9010 16590 9100 16830
rect 9340 16590 9430 16830
rect 9670 16590 9760 16830
rect 10000 16590 10090 16830
rect 10330 16590 10420 16830
rect 10660 16590 10750 16830
rect 10990 16590 11080 16830
rect 11320 16590 11410 16830
rect 11650 16590 11740 16830
rect 11980 16590 12070 16830
rect 12310 16590 12400 16830
rect 12640 16590 12730 16830
rect 12970 16590 13060 16830
rect 13300 16590 13390 16830
rect 13630 16590 13720 16830
rect 13960 16590 14050 16830
rect 14290 16590 14380 16830
rect 14620 16590 14710 16830
rect 14950 16590 15040 16830
rect 15280 16590 15370 16830
rect 15610 16590 15700 16830
rect 15940 16590 16030 16830
rect 16270 16590 16360 16830
rect 16600 16590 16690 16830
rect 16930 16590 17020 16830
rect 17260 16590 17350 16830
rect 17590 16590 17680 16830
rect 17920 16590 18010 16830
rect 18250 16590 18340 16830
rect 18580 16590 18670 16830
rect 18910 16590 19000 16830
rect 19240 16590 19330 16830
rect 19570 16590 19880 16830
rect 7640 16500 19880 16590
rect 7640 16260 7780 16500
rect 8020 16260 8110 16500
rect 8350 16260 8440 16500
rect 8680 16260 8770 16500
rect 9010 16260 9100 16500
rect 9340 16260 9430 16500
rect 9670 16260 9760 16500
rect 10000 16260 10090 16500
rect 10330 16260 10420 16500
rect 10660 16260 10750 16500
rect 10990 16260 11080 16500
rect 11320 16260 11410 16500
rect 11650 16260 11740 16500
rect 11980 16260 12070 16500
rect 12310 16260 12400 16500
rect 12640 16260 12730 16500
rect 12970 16260 13060 16500
rect 13300 16260 13390 16500
rect 13630 16260 13720 16500
rect 13960 16260 14050 16500
rect 14290 16260 14380 16500
rect 14620 16260 14710 16500
rect 14950 16260 15040 16500
rect 15280 16260 15370 16500
rect 15610 16260 15700 16500
rect 15940 16260 16030 16500
rect 16270 16260 16360 16500
rect 16600 16260 16690 16500
rect 16930 16260 17020 16500
rect 17260 16260 17350 16500
rect 17590 16260 17680 16500
rect 17920 16260 18010 16500
rect 18250 16260 18340 16500
rect 18580 16260 18670 16500
rect 18910 16260 19000 16500
rect 19240 16260 19330 16500
rect 19570 16260 19880 16500
rect 7640 16170 19880 16260
rect 7640 15930 7780 16170
rect 8020 15930 8110 16170
rect 8350 15930 8440 16170
rect 8680 15930 8770 16170
rect 9010 15930 9100 16170
rect 9340 15930 9430 16170
rect 9670 15930 9760 16170
rect 10000 15930 10090 16170
rect 10330 15930 10420 16170
rect 10660 15930 10750 16170
rect 10990 15930 11080 16170
rect 11320 15930 11410 16170
rect 11650 15930 11740 16170
rect 11980 15930 12070 16170
rect 12310 15930 12400 16170
rect 12640 15930 12730 16170
rect 12970 15930 13060 16170
rect 13300 15930 13390 16170
rect 13630 15930 13720 16170
rect 13960 15930 14050 16170
rect 14290 15930 14380 16170
rect 14620 15930 14710 16170
rect 14950 15930 15040 16170
rect 15280 15930 15370 16170
rect 15610 15930 15700 16170
rect 15940 15930 16030 16170
rect 16270 15930 16360 16170
rect 16600 15930 16690 16170
rect 16930 15930 17020 16170
rect 17260 15930 17350 16170
rect 17590 15930 17680 16170
rect 17920 15930 18010 16170
rect 18250 15930 18340 16170
rect 18580 15930 18670 16170
rect 18910 15930 19000 16170
rect 19240 15930 19330 16170
rect 19570 15930 19880 16170
rect 7640 15840 19880 15930
rect 7640 15600 7780 15840
rect 8020 15600 8110 15840
rect 8350 15600 8440 15840
rect 8680 15600 8770 15840
rect 9010 15600 9100 15840
rect 9340 15600 9430 15840
rect 9670 15600 9760 15840
rect 10000 15600 10090 15840
rect 10330 15600 10420 15840
rect 10660 15600 10750 15840
rect 10990 15600 11080 15840
rect 11320 15600 11410 15840
rect 11650 15600 11740 15840
rect 11980 15600 12070 15840
rect 12310 15600 12400 15840
rect 12640 15600 12730 15840
rect 12970 15600 13060 15840
rect 13300 15600 13390 15840
rect 13630 15600 13720 15840
rect 13960 15600 14050 15840
rect 14290 15600 14380 15840
rect 14620 15600 14710 15840
rect 14950 15600 15040 15840
rect 15280 15600 15370 15840
rect 15610 15600 15700 15840
rect 15940 15600 16030 15840
rect 16270 15600 16360 15840
rect 16600 15600 16690 15840
rect 16930 15600 17020 15840
rect 17260 15600 17350 15840
rect 17590 15600 17680 15840
rect 17920 15600 18010 15840
rect 18250 15600 18340 15840
rect 18580 15600 18670 15840
rect 18910 15600 19000 15840
rect 19240 15600 19330 15840
rect 19570 15600 19880 15840
rect 7640 15510 19880 15600
rect 7640 15270 7780 15510
rect 8020 15270 8110 15510
rect 8350 15270 8440 15510
rect 8680 15270 8770 15510
rect 9010 15270 9100 15510
rect 9340 15270 9430 15510
rect 9670 15270 9760 15510
rect 10000 15270 10090 15510
rect 10330 15270 10420 15510
rect 10660 15270 10750 15510
rect 10990 15270 11080 15510
rect 11320 15270 11410 15510
rect 11650 15270 11740 15510
rect 11980 15270 12070 15510
rect 12310 15270 12400 15510
rect 12640 15270 12730 15510
rect 12970 15270 13060 15510
rect 13300 15270 13390 15510
rect 13630 15270 13720 15510
rect 13960 15270 14050 15510
rect 14290 15270 14380 15510
rect 14620 15270 14710 15510
rect 14950 15270 15040 15510
rect 15280 15270 15370 15510
rect 15610 15270 15700 15510
rect 15940 15270 16030 15510
rect 16270 15270 16360 15510
rect 16600 15270 16690 15510
rect 16930 15270 17020 15510
rect 17260 15270 17350 15510
rect 17590 15270 17680 15510
rect 17920 15270 18010 15510
rect 18250 15270 18340 15510
rect 18580 15270 18670 15510
rect 18910 15270 19000 15510
rect 19240 15270 19330 15510
rect 19570 15270 19880 15510
rect 7640 15180 19880 15270
rect 7640 14940 7780 15180
rect 8020 14940 8110 15180
rect 8350 14940 8440 15180
rect 8680 14940 8770 15180
rect 9010 14940 9100 15180
rect 9340 14940 9430 15180
rect 9670 14940 9760 15180
rect 10000 14940 10090 15180
rect 10330 14940 10420 15180
rect 10660 14940 10750 15180
rect 10990 14940 11080 15180
rect 11320 14940 11410 15180
rect 11650 14940 11740 15180
rect 11980 14940 12070 15180
rect 12310 14940 12400 15180
rect 12640 14940 12730 15180
rect 12970 14940 13060 15180
rect 13300 14940 13390 15180
rect 13630 14940 13720 15180
rect 13960 14940 14050 15180
rect 14290 14940 14380 15180
rect 14620 14940 14710 15180
rect 14950 14940 15040 15180
rect 15280 14940 15370 15180
rect 15610 14940 15700 15180
rect 15940 14940 16030 15180
rect 16270 14940 16360 15180
rect 16600 14940 16690 15180
rect 16930 14940 17020 15180
rect 17260 14940 17350 15180
rect 17590 14940 17680 15180
rect 17920 14940 18010 15180
rect 18250 14940 18340 15180
rect 18580 14940 18670 15180
rect 18910 14940 19000 15180
rect 19240 14940 19330 15180
rect 19570 14940 19880 15180
rect 7640 14850 19880 14940
rect 7640 14610 7780 14850
rect 8020 14610 8110 14850
rect 8350 14610 8440 14850
rect 8680 14610 8770 14850
rect 9010 14610 9100 14850
rect 9340 14610 9430 14850
rect 9670 14610 9760 14850
rect 10000 14610 10090 14850
rect 10330 14610 10420 14850
rect 10660 14610 10750 14850
rect 10990 14610 11080 14850
rect 11320 14610 11410 14850
rect 11650 14610 11740 14850
rect 11980 14610 12070 14850
rect 12310 14610 12400 14850
rect 12640 14610 12730 14850
rect 12970 14610 13060 14850
rect 13300 14610 13390 14850
rect 13630 14610 13720 14850
rect 13960 14610 14050 14850
rect 14290 14610 14380 14850
rect 14620 14610 14710 14850
rect 14950 14610 15040 14850
rect 15280 14610 15370 14850
rect 15610 14610 15700 14850
rect 15940 14610 16030 14850
rect 16270 14610 16360 14850
rect 16600 14610 16690 14850
rect 16930 14610 17020 14850
rect 17260 14610 17350 14850
rect 17590 14610 17680 14850
rect 17920 14610 18010 14850
rect 18250 14610 18340 14850
rect 18580 14610 18670 14850
rect 18910 14610 19000 14850
rect 19240 14610 19330 14850
rect 19570 14610 19880 14850
rect 7640 14520 19880 14610
rect 7640 14280 7780 14520
rect 8020 14280 8110 14520
rect 8350 14280 8440 14520
rect 8680 14280 8770 14520
rect 9010 14280 9100 14520
rect 9340 14280 9430 14520
rect 9670 14280 9760 14520
rect 10000 14280 10090 14520
rect 10330 14280 10420 14520
rect 10660 14280 10750 14520
rect 10990 14280 11080 14520
rect 11320 14280 11410 14520
rect 11650 14280 11740 14520
rect 11980 14280 12070 14520
rect 12310 14280 12400 14520
rect 12640 14280 12730 14520
rect 12970 14280 13060 14520
rect 13300 14280 13390 14520
rect 13630 14280 13720 14520
rect 13960 14280 14050 14520
rect 14290 14280 14380 14520
rect 14620 14280 14710 14520
rect 14950 14280 15040 14520
rect 15280 14280 15370 14520
rect 15610 14280 15700 14520
rect 15940 14280 16030 14520
rect 16270 14280 16360 14520
rect 16600 14280 16690 14520
rect 16930 14280 17020 14520
rect 17260 14280 17350 14520
rect 17590 14280 17680 14520
rect 17920 14280 18010 14520
rect 18250 14280 18340 14520
rect 18580 14280 18670 14520
rect 18910 14280 19000 14520
rect 19240 14280 19330 14520
rect 19570 14280 19880 14520
rect 7640 14190 19880 14280
rect 7640 13950 7780 14190
rect 8020 13950 8110 14190
rect 8350 13950 8440 14190
rect 8680 13950 8770 14190
rect 9010 13950 9100 14190
rect 9340 13950 9430 14190
rect 9670 13950 9760 14190
rect 10000 13950 10090 14190
rect 10330 13950 10420 14190
rect 10660 13950 10750 14190
rect 10990 13950 11080 14190
rect 11320 13950 11410 14190
rect 11650 13950 11740 14190
rect 11980 13950 12070 14190
rect 12310 13950 12400 14190
rect 12640 13950 12730 14190
rect 12970 13950 13060 14190
rect 13300 13950 13390 14190
rect 13630 13950 13720 14190
rect 13960 13950 14050 14190
rect 14290 13950 14380 14190
rect 14620 13950 14710 14190
rect 14950 13950 15040 14190
rect 15280 13950 15370 14190
rect 15610 13950 15700 14190
rect 15940 13950 16030 14190
rect 16270 13950 16360 14190
rect 16600 13950 16690 14190
rect 16930 13950 17020 14190
rect 17260 13950 17350 14190
rect 17590 13950 17680 14190
rect 17920 13950 18010 14190
rect 18250 13950 18340 14190
rect 18580 13950 18670 14190
rect 18910 13950 19000 14190
rect 19240 13950 19330 14190
rect 19570 13950 19880 14190
rect 7640 13860 19880 13950
rect 7640 13620 7780 13860
rect 8020 13620 8110 13860
rect 8350 13620 8440 13860
rect 8680 13620 8770 13860
rect 9010 13620 9100 13860
rect 9340 13620 9430 13860
rect 9670 13620 9760 13860
rect 10000 13620 10090 13860
rect 10330 13620 10420 13860
rect 10660 13620 10750 13860
rect 10990 13620 11080 13860
rect 11320 13620 11410 13860
rect 11650 13620 11740 13860
rect 11980 13620 12070 13860
rect 12310 13620 12400 13860
rect 12640 13620 12730 13860
rect 12970 13620 13060 13860
rect 13300 13620 13390 13860
rect 13630 13620 13720 13860
rect 13960 13620 14050 13860
rect 14290 13620 14380 13860
rect 14620 13620 14710 13860
rect 14950 13620 15040 13860
rect 15280 13620 15370 13860
rect 15610 13620 15700 13860
rect 15940 13620 16030 13860
rect 16270 13620 16360 13860
rect 16600 13620 16690 13860
rect 16930 13620 17020 13860
rect 17260 13620 17350 13860
rect 17590 13620 17680 13860
rect 17920 13620 18010 13860
rect 18250 13620 18340 13860
rect 18580 13620 18670 13860
rect 18910 13620 19000 13860
rect 19240 13620 19330 13860
rect 19570 13620 19880 13860
rect 7640 13530 19880 13620
rect 7640 13290 7780 13530
rect 8020 13290 8110 13530
rect 8350 13290 8440 13530
rect 8680 13290 8770 13530
rect 9010 13290 9100 13530
rect 9340 13290 9430 13530
rect 9670 13290 9760 13530
rect 10000 13290 10090 13530
rect 10330 13290 10420 13530
rect 10660 13290 10750 13530
rect 10990 13290 11080 13530
rect 11320 13290 11410 13530
rect 11650 13290 11740 13530
rect 11980 13290 12070 13530
rect 12310 13290 12400 13530
rect 12640 13290 12730 13530
rect 12970 13290 13060 13530
rect 13300 13290 13390 13530
rect 13630 13290 13720 13530
rect 13960 13290 14050 13530
rect 14290 13290 14380 13530
rect 14620 13290 14710 13530
rect 14950 13290 15040 13530
rect 15280 13290 15370 13530
rect 15610 13290 15700 13530
rect 15940 13290 16030 13530
rect 16270 13290 16360 13530
rect 16600 13290 16690 13530
rect 16930 13290 17020 13530
rect 17260 13290 17350 13530
rect 17590 13290 17680 13530
rect 17920 13290 18010 13530
rect 18250 13290 18340 13530
rect 18580 13290 18670 13530
rect 18910 13290 19000 13530
rect 19240 13290 19330 13530
rect 19570 13290 19880 13530
rect 7640 13200 19880 13290
rect 7640 12960 7780 13200
rect 8020 12960 8110 13200
rect 8350 12960 8440 13200
rect 8680 12960 8770 13200
rect 9010 12960 9100 13200
rect 9340 12960 9430 13200
rect 9670 12960 9760 13200
rect 10000 12960 10090 13200
rect 10330 12960 10420 13200
rect 10660 12960 10750 13200
rect 10990 12960 11080 13200
rect 11320 12960 11410 13200
rect 11650 12960 11740 13200
rect 11980 12960 12070 13200
rect 12310 12960 12400 13200
rect 12640 12960 12730 13200
rect 12970 12960 13060 13200
rect 13300 12960 13390 13200
rect 13630 12960 13720 13200
rect 13960 12960 14050 13200
rect 14290 12960 14380 13200
rect 14620 12960 14710 13200
rect 14950 12960 15040 13200
rect 15280 12960 15370 13200
rect 15610 12960 15700 13200
rect 15940 12960 16030 13200
rect 16270 12960 16360 13200
rect 16600 12960 16690 13200
rect 16930 12960 17020 13200
rect 17260 12960 17350 13200
rect 17590 12960 17680 13200
rect 17920 12960 18010 13200
rect 18250 12960 18340 13200
rect 18580 12960 18670 13200
rect 18910 12960 19000 13200
rect 19240 12960 19330 13200
rect 19570 12960 19880 13200
rect 7640 12870 19880 12960
rect 7640 12630 7780 12870
rect 8020 12630 8110 12870
rect 8350 12630 8440 12870
rect 8680 12630 8770 12870
rect 9010 12630 9100 12870
rect 9340 12630 9430 12870
rect 9670 12630 9760 12870
rect 10000 12630 10090 12870
rect 10330 12630 10420 12870
rect 10660 12630 10750 12870
rect 10990 12630 11080 12870
rect 11320 12630 11410 12870
rect 11650 12630 11740 12870
rect 11980 12630 12070 12870
rect 12310 12630 12400 12870
rect 12640 12630 12730 12870
rect 12970 12630 13060 12870
rect 13300 12630 13390 12870
rect 13630 12630 13720 12870
rect 13960 12630 14050 12870
rect 14290 12630 14380 12870
rect 14620 12630 14710 12870
rect 14950 12630 15040 12870
rect 15280 12630 15370 12870
rect 15610 12630 15700 12870
rect 15940 12630 16030 12870
rect 16270 12630 16360 12870
rect 16600 12630 16690 12870
rect 16930 12630 17020 12870
rect 17260 12630 17350 12870
rect 17590 12630 17680 12870
rect 17920 12630 18010 12870
rect 18250 12630 18340 12870
rect 18580 12630 18670 12870
rect 18910 12630 19000 12870
rect 19240 12630 19330 12870
rect 19570 12630 19880 12870
rect 7640 12540 19880 12630
rect 7640 12300 7780 12540
rect 8020 12300 8110 12540
rect 8350 12300 8440 12540
rect 8680 12300 8770 12540
rect 9010 12300 9100 12540
rect 9340 12300 9430 12540
rect 9670 12300 9760 12540
rect 10000 12300 10090 12540
rect 10330 12300 10420 12540
rect 10660 12300 10750 12540
rect 10990 12300 11080 12540
rect 11320 12300 11410 12540
rect 11650 12300 11740 12540
rect 11980 12300 12070 12540
rect 12310 12300 12400 12540
rect 12640 12300 12730 12540
rect 12970 12300 13060 12540
rect 13300 12300 13390 12540
rect 13630 12300 13720 12540
rect 13960 12300 14050 12540
rect 14290 12300 14380 12540
rect 14620 12300 14710 12540
rect 14950 12300 15040 12540
rect 15280 12300 15370 12540
rect 15610 12300 15700 12540
rect 15940 12300 16030 12540
rect 16270 12300 16360 12540
rect 16600 12300 16690 12540
rect 16930 12300 17020 12540
rect 17260 12300 17350 12540
rect 17590 12300 17680 12540
rect 17920 12300 18010 12540
rect 18250 12300 18340 12540
rect 18580 12300 18670 12540
rect 18910 12300 19000 12540
rect 19240 12300 19330 12540
rect 19570 12300 19880 12540
rect 7640 12210 19880 12300
rect 7640 11970 7780 12210
rect 8020 11970 8110 12210
rect 8350 11970 8440 12210
rect 8680 11970 8770 12210
rect 9010 11970 9100 12210
rect 9340 11970 9430 12210
rect 9670 11970 9760 12210
rect 10000 11970 10090 12210
rect 10330 11970 10420 12210
rect 10660 11970 10750 12210
rect 10990 11970 11080 12210
rect 11320 11970 11410 12210
rect 11650 11970 11740 12210
rect 11980 11970 12070 12210
rect 12310 11970 12400 12210
rect 12640 11970 12730 12210
rect 12970 11970 13060 12210
rect 13300 11970 13390 12210
rect 13630 11970 13720 12210
rect 13960 11970 14050 12210
rect 14290 11970 14380 12210
rect 14620 11970 14710 12210
rect 14950 11970 15040 12210
rect 15280 11970 15370 12210
rect 15610 11970 15700 12210
rect 15940 11970 16030 12210
rect 16270 11970 16360 12210
rect 16600 11970 16690 12210
rect 16930 11970 17020 12210
rect 17260 11970 17350 12210
rect 17590 11970 17680 12210
rect 17920 11970 18010 12210
rect 18250 11970 18340 12210
rect 18580 11970 18670 12210
rect 18910 11970 19000 12210
rect 19240 11970 19330 12210
rect 19570 11970 19880 12210
rect 7640 11880 19880 11970
rect 7640 11640 7780 11880
rect 8020 11640 8110 11880
rect 8350 11640 8440 11880
rect 8680 11640 8770 11880
rect 9010 11640 9100 11880
rect 9340 11640 9430 11880
rect 9670 11640 9760 11880
rect 10000 11640 10090 11880
rect 10330 11640 10420 11880
rect 10660 11640 10750 11880
rect 10990 11640 11080 11880
rect 11320 11640 11410 11880
rect 11650 11640 11740 11880
rect 11980 11640 12070 11880
rect 12310 11640 12400 11880
rect 12640 11640 12730 11880
rect 12970 11640 13060 11880
rect 13300 11640 13390 11880
rect 13630 11640 13720 11880
rect 13960 11640 14050 11880
rect 14290 11640 14380 11880
rect 14620 11640 14710 11880
rect 14950 11640 15040 11880
rect 15280 11640 15370 11880
rect 15610 11640 15700 11880
rect 15940 11640 16030 11880
rect 16270 11640 16360 11880
rect 16600 11640 16690 11880
rect 16930 11640 17020 11880
rect 17260 11640 17350 11880
rect 17590 11640 17680 11880
rect 17920 11640 18010 11880
rect 18250 11640 18340 11880
rect 18580 11640 18670 11880
rect 18910 11640 19000 11880
rect 19240 11640 19330 11880
rect 19570 11640 19880 11880
rect 7640 11550 19880 11640
rect 7640 11310 7780 11550
rect 8020 11310 8110 11550
rect 8350 11310 8440 11550
rect 8680 11310 8770 11550
rect 9010 11310 9100 11550
rect 9340 11310 9430 11550
rect 9670 11310 9760 11550
rect 10000 11310 10090 11550
rect 10330 11310 10420 11550
rect 10660 11310 10750 11550
rect 10990 11310 11080 11550
rect 11320 11310 11410 11550
rect 11650 11310 11740 11550
rect 11980 11310 12070 11550
rect 12310 11310 12400 11550
rect 12640 11310 12730 11550
rect 12970 11310 13060 11550
rect 13300 11310 13390 11550
rect 13630 11310 13720 11550
rect 13960 11310 14050 11550
rect 14290 11310 14380 11550
rect 14620 11310 14710 11550
rect 14950 11310 15040 11550
rect 15280 11310 15370 11550
rect 15610 11310 15700 11550
rect 15940 11310 16030 11550
rect 16270 11310 16360 11550
rect 16600 11310 16690 11550
rect 16930 11310 17020 11550
rect 17260 11310 17350 11550
rect 17590 11310 17680 11550
rect 17920 11310 18010 11550
rect 18250 11310 18340 11550
rect 18580 11310 18670 11550
rect 18910 11310 19000 11550
rect 19240 11310 19330 11550
rect 19570 11310 19880 11550
rect 7640 11220 19880 11310
rect 7640 10980 7780 11220
rect 8020 10980 8110 11220
rect 8350 10980 8440 11220
rect 8680 10980 8770 11220
rect 9010 10980 9100 11220
rect 9340 10980 9430 11220
rect 9670 10980 9760 11220
rect 10000 10980 10090 11220
rect 10330 10980 10420 11220
rect 10660 10980 10750 11220
rect 10990 10980 11080 11220
rect 11320 10980 11410 11220
rect 11650 10980 11740 11220
rect 11980 10980 12070 11220
rect 12310 10980 12400 11220
rect 12640 10980 12730 11220
rect 12970 10980 13060 11220
rect 13300 10980 13390 11220
rect 13630 10980 13720 11220
rect 13960 10980 14050 11220
rect 14290 10980 14380 11220
rect 14620 10980 14710 11220
rect 14950 10980 15040 11220
rect 15280 10980 15370 11220
rect 15610 10980 15700 11220
rect 15940 10980 16030 11220
rect 16270 10980 16360 11220
rect 16600 10980 16690 11220
rect 16930 10980 17020 11220
rect 17260 10980 17350 11220
rect 17590 10980 17680 11220
rect 17920 10980 18010 11220
rect 18250 10980 18340 11220
rect 18580 10980 18670 11220
rect 18910 10980 19000 11220
rect 19240 10980 19330 11220
rect 19570 10980 19880 11220
rect 7640 10890 19880 10980
rect 7640 10650 7780 10890
rect 8020 10650 8110 10890
rect 8350 10650 8440 10890
rect 8680 10650 8770 10890
rect 9010 10650 9100 10890
rect 9340 10650 9430 10890
rect 9670 10650 9760 10890
rect 10000 10650 10090 10890
rect 10330 10650 10420 10890
rect 10660 10650 10750 10890
rect 10990 10650 11080 10890
rect 11320 10650 11410 10890
rect 11650 10650 11740 10890
rect 11980 10650 12070 10890
rect 12310 10650 12400 10890
rect 12640 10650 12730 10890
rect 12970 10650 13060 10890
rect 13300 10650 13390 10890
rect 13630 10650 13720 10890
rect 13960 10650 14050 10890
rect 14290 10650 14380 10890
rect 14620 10650 14710 10890
rect 14950 10650 15040 10890
rect 15280 10650 15370 10890
rect 15610 10650 15700 10890
rect 15940 10650 16030 10890
rect 16270 10650 16360 10890
rect 16600 10650 16690 10890
rect 16930 10650 17020 10890
rect 17260 10650 17350 10890
rect 17590 10650 17680 10890
rect 17920 10650 18010 10890
rect 18250 10650 18340 10890
rect 18580 10650 18670 10890
rect 18910 10650 19000 10890
rect 19240 10650 19330 10890
rect 19570 10650 19880 10890
rect 7640 10560 19880 10650
rect 7640 10320 7780 10560
rect 8020 10320 8110 10560
rect 8350 10320 8440 10560
rect 8680 10320 8770 10560
rect 9010 10320 9100 10560
rect 9340 10320 9430 10560
rect 9670 10320 9760 10560
rect 10000 10320 10090 10560
rect 10330 10320 10420 10560
rect 10660 10320 10750 10560
rect 10990 10320 11080 10560
rect 11320 10320 11410 10560
rect 11650 10320 11740 10560
rect 11980 10320 12070 10560
rect 12310 10320 12400 10560
rect 12640 10320 12730 10560
rect 12970 10320 13060 10560
rect 13300 10320 13390 10560
rect 13630 10320 13720 10560
rect 13960 10320 14050 10560
rect 14290 10320 14380 10560
rect 14620 10320 14710 10560
rect 14950 10320 15040 10560
rect 15280 10320 15370 10560
rect 15610 10320 15700 10560
rect 15940 10320 16030 10560
rect 16270 10320 16360 10560
rect 16600 10320 16690 10560
rect 16930 10320 17020 10560
rect 17260 10320 17350 10560
rect 17590 10320 17680 10560
rect 17920 10320 18010 10560
rect 18250 10320 18340 10560
rect 18580 10320 18670 10560
rect 18910 10320 19000 10560
rect 19240 10320 19330 10560
rect 19570 10320 19880 10560
rect 7640 10230 19880 10320
rect 7640 9990 7780 10230
rect 8020 9990 8110 10230
rect 8350 9990 8440 10230
rect 8680 9990 8770 10230
rect 9010 9990 9100 10230
rect 9340 9990 9430 10230
rect 9670 9990 9760 10230
rect 10000 9990 10090 10230
rect 10330 9990 10420 10230
rect 10660 9990 10750 10230
rect 10990 9990 11080 10230
rect 11320 9990 11410 10230
rect 11650 9990 11740 10230
rect 11980 9990 12070 10230
rect 12310 9990 12400 10230
rect 12640 9990 12730 10230
rect 12970 9990 13060 10230
rect 13300 9990 13390 10230
rect 13630 9990 13720 10230
rect 13960 9990 14050 10230
rect 14290 9990 14380 10230
rect 14620 9990 14710 10230
rect 14950 9990 15040 10230
rect 15280 9990 15370 10230
rect 15610 9990 15700 10230
rect 15940 9990 16030 10230
rect 16270 9990 16360 10230
rect 16600 9990 16690 10230
rect 16930 9990 17020 10230
rect 17260 9990 17350 10230
rect 17590 9990 17680 10230
rect 17920 9990 18010 10230
rect 18250 9990 18340 10230
rect 18580 9990 18670 10230
rect 18910 9990 19000 10230
rect 19240 9990 19330 10230
rect 19570 9990 19880 10230
rect 7640 9900 19880 9990
rect 7640 9660 7780 9900
rect 8020 9660 8110 9900
rect 8350 9660 8440 9900
rect 8680 9660 8770 9900
rect 9010 9660 9100 9900
rect 9340 9660 9430 9900
rect 9670 9660 9760 9900
rect 10000 9660 10090 9900
rect 10330 9660 10420 9900
rect 10660 9660 10750 9900
rect 10990 9660 11080 9900
rect 11320 9660 11410 9900
rect 11650 9660 11740 9900
rect 11980 9660 12070 9900
rect 12310 9660 12400 9900
rect 12640 9660 12730 9900
rect 12970 9660 13060 9900
rect 13300 9660 13390 9900
rect 13630 9660 13720 9900
rect 13960 9660 14050 9900
rect 14290 9660 14380 9900
rect 14620 9660 14710 9900
rect 14950 9660 15040 9900
rect 15280 9660 15370 9900
rect 15610 9660 15700 9900
rect 15940 9660 16030 9900
rect 16270 9660 16360 9900
rect 16600 9660 16690 9900
rect 16930 9660 17020 9900
rect 17260 9660 17350 9900
rect 17590 9660 17680 9900
rect 17920 9660 18010 9900
rect 18250 9660 18340 9900
rect 18580 9660 18670 9900
rect 18910 9660 19000 9900
rect 19240 9660 19330 9900
rect 19570 9660 19880 9900
rect 7640 9570 19880 9660
rect 7640 9330 7780 9570
rect 8020 9330 8110 9570
rect 8350 9330 8440 9570
rect 8680 9330 8770 9570
rect 9010 9330 9100 9570
rect 9340 9330 9430 9570
rect 9670 9330 9760 9570
rect 10000 9330 10090 9570
rect 10330 9330 10420 9570
rect 10660 9330 10750 9570
rect 10990 9330 11080 9570
rect 11320 9330 11410 9570
rect 11650 9330 11740 9570
rect 11980 9330 12070 9570
rect 12310 9330 12400 9570
rect 12640 9330 12730 9570
rect 12970 9330 13060 9570
rect 13300 9330 13390 9570
rect 13630 9330 13720 9570
rect 13960 9330 14050 9570
rect 14290 9330 14380 9570
rect 14620 9330 14710 9570
rect 14950 9330 15040 9570
rect 15280 9330 15370 9570
rect 15610 9330 15700 9570
rect 15940 9330 16030 9570
rect 16270 9330 16360 9570
rect 16600 9330 16690 9570
rect 16930 9330 17020 9570
rect 17260 9330 17350 9570
rect 17590 9330 17680 9570
rect 17920 9330 18010 9570
rect 18250 9330 18340 9570
rect 18580 9330 18670 9570
rect 18910 9330 19000 9570
rect 19240 9330 19330 9570
rect 19570 9330 19880 9570
rect 7640 9240 19880 9330
rect 7640 9000 7780 9240
rect 8020 9000 8110 9240
rect 8350 9000 8440 9240
rect 8680 9000 8770 9240
rect 9010 9000 9100 9240
rect 9340 9000 9430 9240
rect 9670 9000 9760 9240
rect 10000 9000 10090 9240
rect 10330 9000 10420 9240
rect 10660 9000 10750 9240
rect 10990 9000 11080 9240
rect 11320 9000 11410 9240
rect 11650 9000 11740 9240
rect 11980 9000 12070 9240
rect 12310 9000 12400 9240
rect 12640 9000 12730 9240
rect 12970 9000 13060 9240
rect 13300 9000 13390 9240
rect 13630 9000 13720 9240
rect 13960 9000 14050 9240
rect 14290 9000 14380 9240
rect 14620 9000 14710 9240
rect 14950 9000 15040 9240
rect 15280 9000 15370 9240
rect 15610 9000 15700 9240
rect 15940 9000 16030 9240
rect 16270 9000 16360 9240
rect 16600 9000 16690 9240
rect 16930 9000 17020 9240
rect 17260 9000 17350 9240
rect 17590 9000 17680 9240
rect 17920 9000 18010 9240
rect 18250 9000 18340 9240
rect 18580 9000 18670 9240
rect 18910 9000 19000 9240
rect 19240 9000 19330 9240
rect 19570 9000 19880 9240
rect 7640 8870 19880 9000
rect 28730 7830 35430 7880
rect 28730 7590 28780 7830
rect 29020 7590 29110 7830
rect 29350 7590 29440 7830
rect 29680 7590 29770 7830
rect 30010 7590 30100 7830
rect 30340 7590 30430 7830
rect 30670 7590 30760 7830
rect 31000 7590 31090 7830
rect 31330 7590 31420 7830
rect 31660 7590 31750 7830
rect 31990 7590 32080 7830
rect 32320 7590 32410 7830
rect 32650 7590 32740 7830
rect 32980 7590 33070 7830
rect 33310 7590 33400 7830
rect 33640 7590 33730 7830
rect 33970 7590 34060 7830
rect 34300 7590 34390 7830
rect 34630 7590 34720 7830
rect 34960 7590 35050 7830
rect 35290 7590 35430 7830
rect 28730 7500 35430 7590
rect 28730 7260 28780 7500
rect 29020 7260 29110 7500
rect 29350 7260 29440 7500
rect 29680 7260 29770 7500
rect 30010 7260 30100 7500
rect 30340 7260 30430 7500
rect 30670 7260 30760 7500
rect 31000 7260 31090 7500
rect 31330 7260 31420 7500
rect 31660 7260 31750 7500
rect 31990 7260 32080 7500
rect 32320 7260 32410 7500
rect 32650 7260 32740 7500
rect 32980 7260 33070 7500
rect 33310 7260 33400 7500
rect 33640 7260 33730 7500
rect 33970 7260 34060 7500
rect 34300 7260 34390 7500
rect 34630 7260 34720 7500
rect 34960 7260 35050 7500
rect 35290 7260 35430 7500
rect 28730 7170 35430 7260
rect 28730 6930 28780 7170
rect 29020 6930 29110 7170
rect 29350 6930 29440 7170
rect 29680 6930 29770 7170
rect 30010 6930 30100 7170
rect 30340 6930 30430 7170
rect 30670 6930 30760 7170
rect 31000 6930 31090 7170
rect 31330 6930 31420 7170
rect 31660 6930 31750 7170
rect 31990 6930 32080 7170
rect 32320 6930 32410 7170
rect 32650 6930 32740 7170
rect 32980 6930 33070 7170
rect 33310 6930 33400 7170
rect 33640 6930 33730 7170
rect 33970 6930 34060 7170
rect 34300 6930 34390 7170
rect 34630 6930 34720 7170
rect 34960 6930 35050 7170
rect 35290 6930 35430 7170
rect 28730 6840 35430 6930
rect 28730 6600 28780 6840
rect 29020 6600 29110 6840
rect 29350 6600 29440 6840
rect 29680 6600 29770 6840
rect 30010 6600 30100 6840
rect 30340 6600 30430 6840
rect 30670 6600 30760 6840
rect 31000 6600 31090 6840
rect 31330 6600 31420 6840
rect 31660 6600 31750 6840
rect 31990 6600 32080 6840
rect 32320 6600 32410 6840
rect 32650 6600 32740 6840
rect 32980 6600 33070 6840
rect 33310 6600 33400 6840
rect 33640 6600 33730 6840
rect 33970 6600 34060 6840
rect 34300 6600 34390 6840
rect 34630 6600 34720 6840
rect 34960 6600 35050 6840
rect 35290 6600 35430 6840
rect 28730 6510 35430 6600
rect 28730 6270 28780 6510
rect 29020 6270 29110 6510
rect 29350 6270 29440 6510
rect 29680 6270 29770 6510
rect 30010 6270 30100 6510
rect 30340 6270 30430 6510
rect 30670 6270 30760 6510
rect 31000 6270 31090 6510
rect 31330 6270 31420 6510
rect 31660 6270 31750 6510
rect 31990 6270 32080 6510
rect 32320 6270 32410 6510
rect 32650 6270 32740 6510
rect 32980 6270 33070 6510
rect 33310 6270 33400 6510
rect 33640 6270 33730 6510
rect 33970 6270 34060 6510
rect 34300 6270 34390 6510
rect 34630 6270 34720 6510
rect 34960 6270 35050 6510
rect 35290 6270 35430 6510
rect 28730 6180 35430 6270
rect 28730 5940 28780 6180
rect 29020 5940 29110 6180
rect 29350 5940 29440 6180
rect 29680 5940 29770 6180
rect 30010 5940 30100 6180
rect 30340 5940 30430 6180
rect 30670 5940 30760 6180
rect 31000 5940 31090 6180
rect 31330 5940 31420 6180
rect 31660 5940 31750 6180
rect 31990 5940 32080 6180
rect 32320 5940 32410 6180
rect 32650 5940 32740 6180
rect 32980 5940 33070 6180
rect 33310 5940 33400 6180
rect 33640 5940 33730 6180
rect 33970 5940 34060 6180
rect 34300 5940 34390 6180
rect 34630 5940 34720 6180
rect 34960 5940 35050 6180
rect 35290 5940 35430 6180
rect 28730 5850 35430 5940
rect 28730 5610 28780 5850
rect 29020 5610 29110 5850
rect 29350 5610 29440 5850
rect 29680 5610 29770 5850
rect 30010 5610 30100 5850
rect 30340 5610 30430 5850
rect 30670 5610 30760 5850
rect 31000 5610 31090 5850
rect 31330 5610 31420 5850
rect 31660 5610 31750 5850
rect 31990 5610 32080 5850
rect 32320 5610 32410 5850
rect 32650 5610 32740 5850
rect 32980 5610 33070 5850
rect 33310 5610 33400 5850
rect 33640 5610 33730 5850
rect 33970 5610 34060 5850
rect 34300 5610 34390 5850
rect 34630 5610 34720 5850
rect 34960 5610 35050 5850
rect 35290 5610 35430 5850
rect 28730 5520 35430 5610
rect 28730 5280 28780 5520
rect 29020 5280 29110 5520
rect 29350 5280 29440 5520
rect 29680 5280 29770 5520
rect 30010 5280 30100 5520
rect 30340 5280 30430 5520
rect 30670 5280 30760 5520
rect 31000 5280 31090 5520
rect 31330 5280 31420 5520
rect 31660 5280 31750 5520
rect 31990 5280 32080 5520
rect 32320 5280 32410 5520
rect 32650 5280 32740 5520
rect 32980 5280 33070 5520
rect 33310 5280 33400 5520
rect 33640 5280 33730 5520
rect 33970 5280 34060 5520
rect 34300 5280 34390 5520
rect 34630 5280 34720 5520
rect 34960 5280 35050 5520
rect 35290 5280 35430 5520
rect 28730 5190 35430 5280
rect 28730 4950 28780 5190
rect 29020 4950 29110 5190
rect 29350 4950 29440 5190
rect 29680 4950 29770 5190
rect 30010 4950 30100 5190
rect 30340 4950 30430 5190
rect 30670 4950 30760 5190
rect 31000 4950 31090 5190
rect 31330 4950 31420 5190
rect 31660 4950 31750 5190
rect 31990 4950 32080 5190
rect 32320 4950 32410 5190
rect 32650 4950 32740 5190
rect 32980 4950 33070 5190
rect 33310 4950 33400 5190
rect 33640 4950 33730 5190
rect 33970 4950 34060 5190
rect 34300 4950 34390 5190
rect 34630 4950 34720 5190
rect 34960 4950 35050 5190
rect 35290 4950 35430 5190
rect 28730 4860 35430 4950
rect 28730 4620 28780 4860
rect 29020 4620 29110 4860
rect 29350 4620 29440 4860
rect 29680 4620 29770 4860
rect 30010 4620 30100 4860
rect 30340 4620 30430 4860
rect 30670 4620 30760 4860
rect 31000 4620 31090 4860
rect 31330 4620 31420 4860
rect 31660 4620 31750 4860
rect 31990 4620 32080 4860
rect 32320 4620 32410 4860
rect 32650 4620 32740 4860
rect 32980 4620 33070 4860
rect 33310 4620 33400 4860
rect 33640 4620 33730 4860
rect 33970 4620 34060 4860
rect 34300 4620 34390 4860
rect 34630 4620 34720 4860
rect 34960 4620 35050 4860
rect 35290 4620 35430 4860
rect 28730 4530 35430 4620
rect 28730 4290 28780 4530
rect 29020 4290 29110 4530
rect 29350 4290 29440 4530
rect 29680 4290 29770 4530
rect 30010 4290 30100 4530
rect 30340 4290 30430 4530
rect 30670 4290 30760 4530
rect 31000 4290 31090 4530
rect 31330 4290 31420 4530
rect 31660 4290 31750 4530
rect 31990 4290 32080 4530
rect 32320 4290 32410 4530
rect 32650 4290 32740 4530
rect 32980 4290 33070 4530
rect 33310 4290 33400 4530
rect 33640 4290 33730 4530
rect 33970 4290 34060 4530
rect 34300 4290 34390 4530
rect 34630 4290 34720 4530
rect 34960 4290 35050 4530
rect 35290 4290 35430 4530
rect 28730 4200 35430 4290
rect 28730 3960 28780 4200
rect 29020 3960 29110 4200
rect 29350 3960 29440 4200
rect 29680 3960 29770 4200
rect 30010 3960 30100 4200
rect 30340 3960 30430 4200
rect 30670 3960 30760 4200
rect 31000 3960 31090 4200
rect 31330 3960 31420 4200
rect 31660 3960 31750 4200
rect 31990 3960 32080 4200
rect 32320 3960 32410 4200
rect 32650 3960 32740 4200
rect 32980 3960 33070 4200
rect 33310 3960 33400 4200
rect 33640 3960 33730 4200
rect 33970 3960 34060 4200
rect 34300 3960 34390 4200
rect 34630 3960 34720 4200
rect 34960 3960 35050 4200
rect 35290 3960 35430 4200
rect 28730 3870 35430 3960
rect 28730 3630 28780 3870
rect 29020 3630 29110 3870
rect 29350 3630 29440 3870
rect 29680 3630 29770 3870
rect 30010 3630 30100 3870
rect 30340 3630 30430 3870
rect 30670 3630 30760 3870
rect 31000 3630 31090 3870
rect 31330 3630 31420 3870
rect 31660 3630 31750 3870
rect 31990 3630 32080 3870
rect 32320 3630 32410 3870
rect 32650 3630 32740 3870
rect 32980 3630 33070 3870
rect 33310 3630 33400 3870
rect 33640 3630 33730 3870
rect 33970 3630 34060 3870
rect 34300 3630 34390 3870
rect 34630 3630 34720 3870
rect 34960 3630 35050 3870
rect 35290 3630 35430 3870
rect 28730 3540 35430 3630
rect 28730 3300 28780 3540
rect 29020 3300 29110 3540
rect 29350 3300 29440 3540
rect 29680 3300 29770 3540
rect 30010 3300 30100 3540
rect 30340 3300 30430 3540
rect 30670 3300 30760 3540
rect 31000 3300 31090 3540
rect 31330 3300 31420 3540
rect 31660 3300 31750 3540
rect 31990 3300 32080 3540
rect 32320 3300 32410 3540
rect 32650 3300 32740 3540
rect 32980 3300 33070 3540
rect 33310 3300 33400 3540
rect 33640 3300 33730 3540
rect 33970 3300 34060 3540
rect 34300 3300 34390 3540
rect 34630 3300 34720 3540
rect 34960 3300 35050 3540
rect 35290 3300 35430 3540
rect 28730 3210 35430 3300
rect 28730 2970 28780 3210
rect 29020 2970 29110 3210
rect 29350 2970 29440 3210
rect 29680 2970 29770 3210
rect 30010 2970 30100 3210
rect 30340 2970 30430 3210
rect 30670 2970 30760 3210
rect 31000 2970 31090 3210
rect 31330 2970 31420 3210
rect 31660 2970 31750 3210
rect 31990 2970 32080 3210
rect 32320 2970 32410 3210
rect 32650 2970 32740 3210
rect 32980 2970 33070 3210
rect 33310 2970 33400 3210
rect 33640 2970 33730 3210
rect 33970 2970 34060 3210
rect 34300 2970 34390 3210
rect 34630 2970 34720 3210
rect 34960 2970 35050 3210
rect 35290 2970 35430 3210
rect 28730 2880 35430 2970
rect 28730 2640 28780 2880
rect 29020 2640 29110 2880
rect 29350 2640 29440 2880
rect 29680 2640 29770 2880
rect 30010 2640 30100 2880
rect 30340 2640 30430 2880
rect 30670 2640 30760 2880
rect 31000 2640 31090 2880
rect 31330 2640 31420 2880
rect 31660 2640 31750 2880
rect 31990 2640 32080 2880
rect 32320 2640 32410 2880
rect 32650 2640 32740 2880
rect 32980 2640 33070 2880
rect 33310 2640 33400 2880
rect 33640 2640 33730 2880
rect 33970 2640 34060 2880
rect 34300 2640 34390 2880
rect 34630 2640 34720 2880
rect 34960 2640 35050 2880
rect 35290 2640 35430 2880
rect 28730 2550 35430 2640
rect 28730 2310 28780 2550
rect 29020 2310 29110 2550
rect 29350 2310 29440 2550
rect 29680 2310 29770 2550
rect 30010 2310 30100 2550
rect 30340 2310 30430 2550
rect 30670 2310 30760 2550
rect 31000 2310 31090 2550
rect 31330 2310 31420 2550
rect 31660 2310 31750 2550
rect 31990 2310 32080 2550
rect 32320 2310 32410 2550
rect 32650 2310 32740 2550
rect 32980 2310 33070 2550
rect 33310 2310 33400 2550
rect 33640 2310 33730 2550
rect 33970 2310 34060 2550
rect 34300 2310 34390 2550
rect 34630 2310 34720 2550
rect 34960 2310 35050 2550
rect 35290 2310 35430 2550
rect 28730 2220 35430 2310
rect 28730 1980 28780 2220
rect 29020 1980 29110 2220
rect 29350 1980 29440 2220
rect 29680 1980 29770 2220
rect 30010 1980 30100 2220
rect 30340 1980 30430 2220
rect 30670 1980 30760 2220
rect 31000 1980 31090 2220
rect 31330 1980 31420 2220
rect 31660 1980 31750 2220
rect 31990 1980 32080 2220
rect 32320 1980 32410 2220
rect 32650 1980 32740 2220
rect 32980 1980 33070 2220
rect 33310 1980 33400 2220
rect 33640 1980 33730 2220
rect 33970 1980 34060 2220
rect 34300 1980 34390 2220
rect 34630 1980 34720 2220
rect 34960 1980 35050 2220
rect 35290 1980 35430 2220
rect 28730 1890 35430 1980
rect 28730 1650 28780 1890
rect 29020 1650 29110 1890
rect 29350 1650 29440 1890
rect 29680 1650 29770 1890
rect 30010 1650 30100 1890
rect 30340 1650 30430 1890
rect 30670 1650 30760 1890
rect 31000 1650 31090 1890
rect 31330 1650 31420 1890
rect 31660 1650 31750 1890
rect 31990 1650 32080 1890
rect 32320 1650 32410 1890
rect 32650 1650 32740 1890
rect 32980 1650 33070 1890
rect 33310 1650 33400 1890
rect 33640 1650 33730 1890
rect 33970 1650 34060 1890
rect 34300 1650 34390 1890
rect 34630 1650 34720 1890
rect 34960 1650 35050 1890
rect 35290 1650 35430 1890
rect 28730 1560 35430 1650
rect 28730 1320 28780 1560
rect 29020 1320 29110 1560
rect 29350 1320 29440 1560
rect 29680 1320 29770 1560
rect 30010 1320 30100 1560
rect 30340 1320 30430 1560
rect 30670 1320 30760 1560
rect 31000 1320 31090 1560
rect 31330 1320 31420 1560
rect 31660 1320 31750 1560
rect 31990 1320 32080 1560
rect 32320 1320 32410 1560
rect 32650 1320 32740 1560
rect 32980 1320 33070 1560
rect 33310 1320 33400 1560
rect 33640 1320 33730 1560
rect 33970 1320 34060 1560
rect 34300 1320 34390 1560
rect 34630 1320 34720 1560
rect 34960 1320 35050 1560
rect 35290 1320 35430 1560
rect 28730 1180 35430 1320
rect 28730 230 35430 280
rect 28730 -10 28780 230
rect 29020 -10 29110 230
rect 29350 -10 29440 230
rect 29680 -10 29770 230
rect 30010 -10 30100 230
rect 30340 -10 30430 230
rect 30670 -10 30760 230
rect 31000 -10 31090 230
rect 31330 -10 31420 230
rect 31660 -10 31750 230
rect 31990 -10 32080 230
rect 32320 -10 32410 230
rect 32650 -10 32740 230
rect 32980 -10 33070 230
rect 33310 -10 33400 230
rect 33640 -10 33730 230
rect 33970 -10 34060 230
rect 34300 -10 34390 230
rect 34630 -10 34720 230
rect 34960 -10 35050 230
rect 35290 -10 35430 230
rect 28730 -100 35430 -10
rect 28730 -340 28780 -100
rect 29020 -340 29110 -100
rect 29350 -340 29440 -100
rect 29680 -340 29770 -100
rect 30010 -340 30100 -100
rect 30340 -340 30430 -100
rect 30670 -340 30760 -100
rect 31000 -340 31090 -100
rect 31330 -340 31420 -100
rect 31660 -340 31750 -100
rect 31990 -340 32080 -100
rect 32320 -340 32410 -100
rect 32650 -340 32740 -100
rect 32980 -340 33070 -100
rect 33310 -340 33400 -100
rect 33640 -340 33730 -100
rect 33970 -340 34060 -100
rect 34300 -340 34390 -100
rect 34630 -340 34720 -100
rect 34960 -340 35050 -100
rect 35290 -340 35430 -100
rect 28730 -430 35430 -340
rect 28730 -670 28780 -430
rect 29020 -670 29110 -430
rect 29350 -670 29440 -430
rect 29680 -670 29770 -430
rect 30010 -670 30100 -430
rect 30340 -670 30430 -430
rect 30670 -670 30760 -430
rect 31000 -670 31090 -430
rect 31330 -670 31420 -430
rect 31660 -670 31750 -430
rect 31990 -670 32080 -430
rect 32320 -670 32410 -430
rect 32650 -670 32740 -430
rect 32980 -670 33070 -430
rect 33310 -670 33400 -430
rect 33640 -670 33730 -430
rect 33970 -670 34060 -430
rect 34300 -670 34390 -430
rect 34630 -670 34720 -430
rect 34960 -670 35050 -430
rect 35290 -670 35430 -430
rect 28730 -760 35430 -670
rect 28730 -1000 28780 -760
rect 29020 -1000 29110 -760
rect 29350 -1000 29440 -760
rect 29680 -1000 29770 -760
rect 30010 -1000 30100 -760
rect 30340 -1000 30430 -760
rect 30670 -1000 30760 -760
rect 31000 -1000 31090 -760
rect 31330 -1000 31420 -760
rect 31660 -1000 31750 -760
rect 31990 -1000 32080 -760
rect 32320 -1000 32410 -760
rect 32650 -1000 32740 -760
rect 32980 -1000 33070 -760
rect 33310 -1000 33400 -760
rect 33640 -1000 33730 -760
rect 33970 -1000 34060 -760
rect 34300 -1000 34390 -760
rect 34630 -1000 34720 -760
rect 34960 -1000 35050 -760
rect 35290 -1000 35430 -760
rect 28730 -1090 35430 -1000
rect 28730 -1330 28780 -1090
rect 29020 -1330 29110 -1090
rect 29350 -1330 29440 -1090
rect 29680 -1330 29770 -1090
rect 30010 -1330 30100 -1090
rect 30340 -1330 30430 -1090
rect 30670 -1330 30760 -1090
rect 31000 -1330 31090 -1090
rect 31330 -1330 31420 -1090
rect 31660 -1330 31750 -1090
rect 31990 -1330 32080 -1090
rect 32320 -1330 32410 -1090
rect 32650 -1330 32740 -1090
rect 32980 -1330 33070 -1090
rect 33310 -1330 33400 -1090
rect 33640 -1330 33730 -1090
rect 33970 -1330 34060 -1090
rect 34300 -1330 34390 -1090
rect 34630 -1330 34720 -1090
rect 34960 -1330 35050 -1090
rect 35290 -1330 35430 -1090
rect 28730 -1420 35430 -1330
rect 28730 -1660 28780 -1420
rect 29020 -1660 29110 -1420
rect 29350 -1660 29440 -1420
rect 29680 -1660 29770 -1420
rect 30010 -1660 30100 -1420
rect 30340 -1660 30430 -1420
rect 30670 -1660 30760 -1420
rect 31000 -1660 31090 -1420
rect 31330 -1660 31420 -1420
rect 31660 -1660 31750 -1420
rect 31990 -1660 32080 -1420
rect 32320 -1660 32410 -1420
rect 32650 -1660 32740 -1420
rect 32980 -1660 33070 -1420
rect 33310 -1660 33400 -1420
rect 33640 -1660 33730 -1420
rect 33970 -1660 34060 -1420
rect 34300 -1660 34390 -1420
rect 34630 -1660 34720 -1420
rect 34960 -1660 35050 -1420
rect 35290 -1660 35430 -1420
rect 28730 -1750 35430 -1660
rect 28730 -1990 28780 -1750
rect 29020 -1990 29110 -1750
rect 29350 -1990 29440 -1750
rect 29680 -1990 29770 -1750
rect 30010 -1990 30100 -1750
rect 30340 -1990 30430 -1750
rect 30670 -1990 30760 -1750
rect 31000 -1990 31090 -1750
rect 31330 -1990 31420 -1750
rect 31660 -1990 31750 -1750
rect 31990 -1990 32080 -1750
rect 32320 -1990 32410 -1750
rect 32650 -1990 32740 -1750
rect 32980 -1990 33070 -1750
rect 33310 -1990 33400 -1750
rect 33640 -1990 33730 -1750
rect 33970 -1990 34060 -1750
rect 34300 -1990 34390 -1750
rect 34630 -1990 34720 -1750
rect 34960 -1990 35050 -1750
rect 35290 -1990 35430 -1750
rect 28730 -2080 35430 -1990
rect 28730 -2320 28780 -2080
rect 29020 -2320 29110 -2080
rect 29350 -2320 29440 -2080
rect 29680 -2320 29770 -2080
rect 30010 -2320 30100 -2080
rect 30340 -2320 30430 -2080
rect 30670 -2320 30760 -2080
rect 31000 -2320 31090 -2080
rect 31330 -2320 31420 -2080
rect 31660 -2320 31750 -2080
rect 31990 -2320 32080 -2080
rect 32320 -2320 32410 -2080
rect 32650 -2320 32740 -2080
rect 32980 -2320 33070 -2080
rect 33310 -2320 33400 -2080
rect 33640 -2320 33730 -2080
rect 33970 -2320 34060 -2080
rect 34300 -2320 34390 -2080
rect 34630 -2320 34720 -2080
rect 34960 -2320 35050 -2080
rect 35290 -2320 35430 -2080
rect 28730 -2410 35430 -2320
rect 28730 -2650 28780 -2410
rect 29020 -2650 29110 -2410
rect 29350 -2650 29440 -2410
rect 29680 -2650 29770 -2410
rect 30010 -2650 30100 -2410
rect 30340 -2650 30430 -2410
rect 30670 -2650 30760 -2410
rect 31000 -2650 31090 -2410
rect 31330 -2650 31420 -2410
rect 31660 -2650 31750 -2410
rect 31990 -2650 32080 -2410
rect 32320 -2650 32410 -2410
rect 32650 -2650 32740 -2410
rect 32980 -2650 33070 -2410
rect 33310 -2650 33400 -2410
rect 33640 -2650 33730 -2410
rect 33970 -2650 34060 -2410
rect 34300 -2650 34390 -2410
rect 34630 -2650 34720 -2410
rect 34960 -2650 35050 -2410
rect 35290 -2650 35430 -2410
rect 28730 -2740 35430 -2650
rect 28730 -2980 28780 -2740
rect 29020 -2980 29110 -2740
rect 29350 -2980 29440 -2740
rect 29680 -2980 29770 -2740
rect 30010 -2980 30100 -2740
rect 30340 -2980 30430 -2740
rect 30670 -2980 30760 -2740
rect 31000 -2980 31090 -2740
rect 31330 -2980 31420 -2740
rect 31660 -2980 31750 -2740
rect 31990 -2980 32080 -2740
rect 32320 -2980 32410 -2740
rect 32650 -2980 32740 -2740
rect 32980 -2980 33070 -2740
rect 33310 -2980 33400 -2740
rect 33640 -2980 33730 -2740
rect 33970 -2980 34060 -2740
rect 34300 -2980 34390 -2740
rect 34630 -2980 34720 -2740
rect 34960 -2980 35050 -2740
rect 35290 -2980 35430 -2740
rect 28730 -3070 35430 -2980
rect 28730 -3310 28780 -3070
rect 29020 -3310 29110 -3070
rect 29350 -3310 29440 -3070
rect 29680 -3310 29770 -3070
rect 30010 -3310 30100 -3070
rect 30340 -3310 30430 -3070
rect 30670 -3310 30760 -3070
rect 31000 -3310 31090 -3070
rect 31330 -3310 31420 -3070
rect 31660 -3310 31750 -3070
rect 31990 -3310 32080 -3070
rect 32320 -3310 32410 -3070
rect 32650 -3310 32740 -3070
rect 32980 -3310 33070 -3070
rect 33310 -3310 33400 -3070
rect 33640 -3310 33730 -3070
rect 33970 -3310 34060 -3070
rect 34300 -3310 34390 -3070
rect 34630 -3310 34720 -3070
rect 34960 -3310 35050 -3070
rect 35290 -3310 35430 -3070
rect 28730 -3400 35430 -3310
rect 28730 -3640 28780 -3400
rect 29020 -3640 29110 -3400
rect 29350 -3640 29440 -3400
rect 29680 -3640 29770 -3400
rect 30010 -3640 30100 -3400
rect 30340 -3640 30430 -3400
rect 30670 -3640 30760 -3400
rect 31000 -3640 31090 -3400
rect 31330 -3640 31420 -3400
rect 31660 -3640 31750 -3400
rect 31990 -3640 32080 -3400
rect 32320 -3640 32410 -3400
rect 32650 -3640 32740 -3400
rect 32980 -3640 33070 -3400
rect 33310 -3640 33400 -3400
rect 33640 -3640 33730 -3400
rect 33970 -3640 34060 -3400
rect 34300 -3640 34390 -3400
rect 34630 -3640 34720 -3400
rect 34960 -3640 35050 -3400
rect 35290 -3640 35430 -3400
rect 28730 -3730 35430 -3640
rect 28730 -3970 28780 -3730
rect 29020 -3970 29110 -3730
rect 29350 -3970 29440 -3730
rect 29680 -3970 29770 -3730
rect 30010 -3970 30100 -3730
rect 30340 -3970 30430 -3730
rect 30670 -3970 30760 -3730
rect 31000 -3970 31090 -3730
rect 31330 -3970 31420 -3730
rect 31660 -3970 31750 -3730
rect 31990 -3970 32080 -3730
rect 32320 -3970 32410 -3730
rect 32650 -3970 32740 -3730
rect 32980 -3970 33070 -3730
rect 33310 -3970 33400 -3730
rect 33640 -3970 33730 -3730
rect 33970 -3970 34060 -3730
rect 34300 -3970 34390 -3730
rect 34630 -3970 34720 -3730
rect 34960 -3970 35050 -3730
rect 35290 -3970 35430 -3730
rect 28730 -4060 35430 -3970
rect -1830 -4260 -280 -4080
rect -1830 -4500 -1650 -4260
rect -1410 -4500 -1320 -4260
rect -1080 -4500 -990 -4260
rect -750 -4500 -660 -4260
rect -420 -4500 -280 -4260
rect -1830 -4590 -280 -4500
rect -1830 -4830 -1650 -4590
rect -1410 -4830 -1320 -4590
rect -1080 -4830 -990 -4590
rect -750 -4830 -660 -4590
rect -420 -4830 -280 -4590
rect -1830 -4920 -280 -4830
rect -1830 -5160 -1650 -4920
rect -1410 -5160 -1320 -4920
rect -1080 -5160 -990 -4920
rect -750 -5160 -660 -4920
rect -420 -5160 -280 -4920
rect -1830 -5250 -280 -5160
rect -1830 -5490 -1650 -5250
rect -1410 -5490 -1320 -5250
rect -1080 -5490 -990 -5250
rect -750 -5490 -660 -5250
rect -420 -5490 -280 -5250
rect -1830 -5630 -280 -5490
rect 28730 -4300 28780 -4060
rect 29020 -4300 29110 -4060
rect 29350 -4300 29440 -4060
rect 29680 -4300 29770 -4060
rect 30010 -4300 30100 -4060
rect 30340 -4300 30430 -4060
rect 30670 -4300 30760 -4060
rect 31000 -4300 31090 -4060
rect 31330 -4300 31420 -4060
rect 31660 -4300 31750 -4060
rect 31990 -4300 32080 -4060
rect 32320 -4300 32410 -4060
rect 32650 -4300 32740 -4060
rect 32980 -4300 33070 -4060
rect 33310 -4300 33400 -4060
rect 33640 -4300 33730 -4060
rect 33970 -4300 34060 -4060
rect 34300 -4300 34390 -4060
rect 34630 -4300 34720 -4060
rect 34960 -4300 35050 -4060
rect 35290 -4300 35430 -4060
rect 28730 -4390 35430 -4300
rect 28730 -4630 28780 -4390
rect 29020 -4630 29110 -4390
rect 29350 -4630 29440 -4390
rect 29680 -4630 29770 -4390
rect 30010 -4630 30100 -4390
rect 30340 -4630 30430 -4390
rect 30670 -4630 30760 -4390
rect 31000 -4630 31090 -4390
rect 31330 -4630 31420 -4390
rect 31660 -4630 31750 -4390
rect 31990 -4630 32080 -4390
rect 32320 -4630 32410 -4390
rect 32650 -4630 32740 -4390
rect 32980 -4630 33070 -4390
rect 33310 -4630 33400 -4390
rect 33640 -4630 33730 -4390
rect 33970 -4630 34060 -4390
rect 34300 -4630 34390 -4390
rect 34630 -4630 34720 -4390
rect 34960 -4630 35050 -4390
rect 35290 -4630 35430 -4390
rect 28730 -4720 35430 -4630
rect 28730 -4960 28780 -4720
rect 29020 -4960 29110 -4720
rect 29350 -4960 29440 -4720
rect 29680 -4960 29770 -4720
rect 30010 -4960 30100 -4720
rect 30340 -4960 30430 -4720
rect 30670 -4960 30760 -4720
rect 31000 -4960 31090 -4720
rect 31330 -4960 31420 -4720
rect 31660 -4960 31750 -4720
rect 31990 -4960 32080 -4720
rect 32320 -4960 32410 -4720
rect 32650 -4960 32740 -4720
rect 32980 -4960 33070 -4720
rect 33310 -4960 33400 -4720
rect 33640 -4960 33730 -4720
rect 33970 -4960 34060 -4720
rect 34300 -4960 34390 -4720
rect 34630 -4960 34720 -4720
rect 34960 -4960 35050 -4720
rect 35290 -4960 35430 -4720
rect 28730 -5050 35430 -4960
rect 28730 -5290 28780 -5050
rect 29020 -5290 29110 -5050
rect 29350 -5290 29440 -5050
rect 29680 -5290 29770 -5050
rect 30010 -5290 30100 -5050
rect 30340 -5290 30430 -5050
rect 30670 -5290 30760 -5050
rect 31000 -5290 31090 -5050
rect 31330 -5290 31420 -5050
rect 31660 -5290 31750 -5050
rect 31990 -5290 32080 -5050
rect 32320 -5290 32410 -5050
rect 32650 -5290 32740 -5050
rect 32980 -5290 33070 -5050
rect 33310 -5290 33400 -5050
rect 33640 -5290 33730 -5050
rect 33970 -5290 34060 -5050
rect 34300 -5290 34390 -5050
rect 34630 -5290 34720 -5050
rect 34960 -5290 35050 -5050
rect 35290 -5290 35430 -5050
rect 28730 -5380 35430 -5290
rect 28730 -5620 28780 -5380
rect 29020 -5620 29110 -5380
rect 29350 -5620 29440 -5380
rect 29680 -5620 29770 -5380
rect 30010 -5620 30100 -5380
rect 30340 -5620 30430 -5380
rect 30670 -5620 30760 -5380
rect 31000 -5620 31090 -5380
rect 31330 -5620 31420 -5380
rect 31660 -5620 31750 -5380
rect 31990 -5620 32080 -5380
rect 32320 -5620 32410 -5380
rect 32650 -5620 32740 -5380
rect 32980 -5620 33070 -5380
rect 33310 -5620 33400 -5380
rect 33640 -5620 33730 -5380
rect 33970 -5620 34060 -5380
rect 34300 -5620 34390 -5380
rect 34630 -5620 34720 -5380
rect 34960 -5620 35050 -5380
rect 35290 -5620 35430 -5380
rect 28730 -5710 35430 -5620
rect 28730 -5950 28780 -5710
rect 29020 -5950 29110 -5710
rect 29350 -5950 29440 -5710
rect 29680 -5950 29770 -5710
rect 30010 -5950 30100 -5710
rect 30340 -5950 30430 -5710
rect 30670 -5950 30760 -5710
rect 31000 -5950 31090 -5710
rect 31330 -5950 31420 -5710
rect 31660 -5950 31750 -5710
rect 31990 -5950 32080 -5710
rect 32320 -5950 32410 -5710
rect 32650 -5950 32740 -5710
rect 32980 -5950 33070 -5710
rect 33310 -5950 33400 -5710
rect 33640 -5950 33730 -5710
rect 33970 -5950 34060 -5710
rect 34300 -5950 34390 -5710
rect 34630 -5950 34720 -5710
rect 34960 -5950 35050 -5710
rect 35290 -5950 35430 -5710
rect 28730 -6040 35430 -5950
rect 28730 -6280 28780 -6040
rect 29020 -6280 29110 -6040
rect 29350 -6280 29440 -6040
rect 29680 -6280 29770 -6040
rect 30010 -6280 30100 -6040
rect 30340 -6280 30430 -6040
rect 30670 -6280 30760 -6040
rect 31000 -6280 31090 -6040
rect 31330 -6280 31420 -6040
rect 31660 -6280 31750 -6040
rect 31990 -6280 32080 -6040
rect 32320 -6280 32410 -6040
rect 32650 -6280 32740 -6040
rect 32980 -6280 33070 -6040
rect 33310 -6280 33400 -6040
rect 33640 -6280 33730 -6040
rect 33970 -6280 34060 -6040
rect 34300 -6280 34390 -6040
rect 34630 -6280 34720 -6040
rect 34960 -6280 35050 -6040
rect 35290 -6280 35430 -6040
rect 28730 -6420 35430 -6280
rect -1830 -7660 -280 -7480
rect -1830 -7900 -1650 -7660
rect -1410 -7900 -1320 -7660
rect -1080 -7900 -990 -7660
rect -750 -7900 -660 -7660
rect -420 -7900 -280 -7660
rect -1830 -7990 -280 -7900
rect -1830 -8230 -1650 -7990
rect -1410 -8230 -1320 -7990
rect -1080 -8230 -990 -7990
rect -750 -8230 -660 -7990
rect -420 -8230 -280 -7990
rect -1830 -8320 -280 -8230
rect -1830 -8560 -1650 -8320
rect -1410 -8560 -1320 -8320
rect -1080 -8560 -990 -8320
rect -750 -8560 -660 -8320
rect -420 -8560 -280 -8320
rect -1830 -8650 -280 -8560
rect -1830 -8890 -1650 -8650
rect -1410 -8890 -1320 -8650
rect -1080 -8890 -990 -8650
rect -750 -8890 -660 -8650
rect -420 -8890 -280 -8650
rect -1830 -9030 -280 -8890
<< mimcapcontact >>
rect -4670 20550 -4430 20790
rect -4340 20550 -4100 20790
rect -4010 20550 -3770 20790
rect -3680 20550 -3440 20790
rect -3350 20550 -3110 20790
rect -3020 20550 -2780 20790
rect -2690 20550 -2450 20790
rect -2360 20550 -2120 20790
rect -2030 20550 -1790 20790
rect -1700 20550 -1460 20790
rect -1370 20550 -1130 20790
rect -1040 20550 -800 20790
rect -710 20550 -470 20790
rect -380 20550 -140 20790
rect -50 20550 190 20790
rect 280 20550 520 20790
rect 610 20550 850 20790
rect 940 20550 1180 20790
rect 1270 20550 1510 20790
rect 1600 20550 1840 20790
rect 1930 20550 2170 20790
rect 2260 20550 2500 20790
rect 2590 20550 2830 20790
rect 2920 20550 3160 20790
rect 3250 20550 3490 20790
rect 3580 20550 3820 20790
rect 3910 20550 4150 20790
rect 4240 20550 4480 20790
rect 4570 20550 4810 20790
rect 4900 20550 5140 20790
rect 5230 20550 5470 20790
rect 5560 20550 5800 20790
rect 5890 20550 6130 20790
rect 6220 20550 6460 20790
rect 6550 20550 6790 20790
rect 6880 20550 7120 20790
rect -4670 20220 -4430 20460
rect -4340 20220 -4100 20460
rect -4010 20220 -3770 20460
rect -3680 20220 -3440 20460
rect -3350 20220 -3110 20460
rect -3020 20220 -2780 20460
rect -2690 20220 -2450 20460
rect -2360 20220 -2120 20460
rect -2030 20220 -1790 20460
rect -1700 20220 -1460 20460
rect -1370 20220 -1130 20460
rect -1040 20220 -800 20460
rect -710 20220 -470 20460
rect -380 20220 -140 20460
rect -50 20220 190 20460
rect 280 20220 520 20460
rect 610 20220 850 20460
rect 940 20220 1180 20460
rect 1270 20220 1510 20460
rect 1600 20220 1840 20460
rect 1930 20220 2170 20460
rect 2260 20220 2500 20460
rect 2590 20220 2830 20460
rect 2920 20220 3160 20460
rect 3250 20220 3490 20460
rect 3580 20220 3820 20460
rect 3910 20220 4150 20460
rect 4240 20220 4480 20460
rect 4570 20220 4810 20460
rect 4900 20220 5140 20460
rect 5230 20220 5470 20460
rect 5560 20220 5800 20460
rect 5890 20220 6130 20460
rect 6220 20220 6460 20460
rect 6550 20220 6790 20460
rect 6880 20220 7120 20460
rect -4670 19890 -4430 20130
rect -4340 19890 -4100 20130
rect -4010 19890 -3770 20130
rect -3680 19890 -3440 20130
rect -3350 19890 -3110 20130
rect -3020 19890 -2780 20130
rect -2690 19890 -2450 20130
rect -2360 19890 -2120 20130
rect -2030 19890 -1790 20130
rect -1700 19890 -1460 20130
rect -1370 19890 -1130 20130
rect -1040 19890 -800 20130
rect -710 19890 -470 20130
rect -380 19890 -140 20130
rect -50 19890 190 20130
rect 280 19890 520 20130
rect 610 19890 850 20130
rect 940 19890 1180 20130
rect 1270 19890 1510 20130
rect 1600 19890 1840 20130
rect 1930 19890 2170 20130
rect 2260 19890 2500 20130
rect 2590 19890 2830 20130
rect 2920 19890 3160 20130
rect 3250 19890 3490 20130
rect 3580 19890 3820 20130
rect 3910 19890 4150 20130
rect 4240 19890 4480 20130
rect 4570 19890 4810 20130
rect 4900 19890 5140 20130
rect 5230 19890 5470 20130
rect 5560 19890 5800 20130
rect 5890 19890 6130 20130
rect 6220 19890 6460 20130
rect 6550 19890 6790 20130
rect 6880 19890 7120 20130
rect -4670 19560 -4430 19800
rect -4340 19560 -4100 19800
rect -4010 19560 -3770 19800
rect -3680 19560 -3440 19800
rect -3350 19560 -3110 19800
rect -3020 19560 -2780 19800
rect -2690 19560 -2450 19800
rect -2360 19560 -2120 19800
rect -2030 19560 -1790 19800
rect -1700 19560 -1460 19800
rect -1370 19560 -1130 19800
rect -1040 19560 -800 19800
rect -710 19560 -470 19800
rect -380 19560 -140 19800
rect -50 19560 190 19800
rect 280 19560 520 19800
rect 610 19560 850 19800
rect 940 19560 1180 19800
rect 1270 19560 1510 19800
rect 1600 19560 1840 19800
rect 1930 19560 2170 19800
rect 2260 19560 2500 19800
rect 2590 19560 2830 19800
rect 2920 19560 3160 19800
rect 3250 19560 3490 19800
rect 3580 19560 3820 19800
rect 3910 19560 4150 19800
rect 4240 19560 4480 19800
rect 4570 19560 4810 19800
rect 4900 19560 5140 19800
rect 5230 19560 5470 19800
rect 5560 19560 5800 19800
rect 5890 19560 6130 19800
rect 6220 19560 6460 19800
rect 6550 19560 6790 19800
rect 6880 19560 7120 19800
rect -4670 19230 -4430 19470
rect -4340 19230 -4100 19470
rect -4010 19230 -3770 19470
rect -3680 19230 -3440 19470
rect -3350 19230 -3110 19470
rect -3020 19230 -2780 19470
rect -2690 19230 -2450 19470
rect -2360 19230 -2120 19470
rect -2030 19230 -1790 19470
rect -1700 19230 -1460 19470
rect -1370 19230 -1130 19470
rect -1040 19230 -800 19470
rect -710 19230 -470 19470
rect -380 19230 -140 19470
rect -50 19230 190 19470
rect 280 19230 520 19470
rect 610 19230 850 19470
rect 940 19230 1180 19470
rect 1270 19230 1510 19470
rect 1600 19230 1840 19470
rect 1930 19230 2170 19470
rect 2260 19230 2500 19470
rect 2590 19230 2830 19470
rect 2920 19230 3160 19470
rect 3250 19230 3490 19470
rect 3580 19230 3820 19470
rect 3910 19230 4150 19470
rect 4240 19230 4480 19470
rect 4570 19230 4810 19470
rect 4900 19230 5140 19470
rect 5230 19230 5470 19470
rect 5560 19230 5800 19470
rect 5890 19230 6130 19470
rect 6220 19230 6460 19470
rect 6550 19230 6790 19470
rect 6880 19230 7120 19470
rect -4670 18900 -4430 19140
rect -4340 18900 -4100 19140
rect -4010 18900 -3770 19140
rect -3680 18900 -3440 19140
rect -3350 18900 -3110 19140
rect -3020 18900 -2780 19140
rect -2690 18900 -2450 19140
rect -2360 18900 -2120 19140
rect -2030 18900 -1790 19140
rect -1700 18900 -1460 19140
rect -1370 18900 -1130 19140
rect -1040 18900 -800 19140
rect -710 18900 -470 19140
rect -380 18900 -140 19140
rect -50 18900 190 19140
rect 280 18900 520 19140
rect 610 18900 850 19140
rect 940 18900 1180 19140
rect 1270 18900 1510 19140
rect 1600 18900 1840 19140
rect 1930 18900 2170 19140
rect 2260 18900 2500 19140
rect 2590 18900 2830 19140
rect 2920 18900 3160 19140
rect 3250 18900 3490 19140
rect 3580 18900 3820 19140
rect 3910 18900 4150 19140
rect 4240 18900 4480 19140
rect 4570 18900 4810 19140
rect 4900 18900 5140 19140
rect 5230 18900 5470 19140
rect 5560 18900 5800 19140
rect 5890 18900 6130 19140
rect 6220 18900 6460 19140
rect 6550 18900 6790 19140
rect 6880 18900 7120 19140
rect -4670 18570 -4430 18810
rect -4340 18570 -4100 18810
rect -4010 18570 -3770 18810
rect -3680 18570 -3440 18810
rect -3350 18570 -3110 18810
rect -3020 18570 -2780 18810
rect -2690 18570 -2450 18810
rect -2360 18570 -2120 18810
rect -2030 18570 -1790 18810
rect -1700 18570 -1460 18810
rect -1370 18570 -1130 18810
rect -1040 18570 -800 18810
rect -710 18570 -470 18810
rect -380 18570 -140 18810
rect -50 18570 190 18810
rect 280 18570 520 18810
rect 610 18570 850 18810
rect 940 18570 1180 18810
rect 1270 18570 1510 18810
rect 1600 18570 1840 18810
rect 1930 18570 2170 18810
rect 2260 18570 2500 18810
rect 2590 18570 2830 18810
rect 2920 18570 3160 18810
rect 3250 18570 3490 18810
rect 3580 18570 3820 18810
rect 3910 18570 4150 18810
rect 4240 18570 4480 18810
rect 4570 18570 4810 18810
rect 4900 18570 5140 18810
rect 5230 18570 5470 18810
rect 5560 18570 5800 18810
rect 5890 18570 6130 18810
rect 6220 18570 6460 18810
rect 6550 18570 6790 18810
rect 6880 18570 7120 18810
rect -4670 18240 -4430 18480
rect -4340 18240 -4100 18480
rect -4010 18240 -3770 18480
rect -3680 18240 -3440 18480
rect -3350 18240 -3110 18480
rect -3020 18240 -2780 18480
rect -2690 18240 -2450 18480
rect -2360 18240 -2120 18480
rect -2030 18240 -1790 18480
rect -1700 18240 -1460 18480
rect -1370 18240 -1130 18480
rect -1040 18240 -800 18480
rect -710 18240 -470 18480
rect -380 18240 -140 18480
rect -50 18240 190 18480
rect 280 18240 520 18480
rect 610 18240 850 18480
rect 940 18240 1180 18480
rect 1270 18240 1510 18480
rect 1600 18240 1840 18480
rect 1930 18240 2170 18480
rect 2260 18240 2500 18480
rect 2590 18240 2830 18480
rect 2920 18240 3160 18480
rect 3250 18240 3490 18480
rect 3580 18240 3820 18480
rect 3910 18240 4150 18480
rect 4240 18240 4480 18480
rect 4570 18240 4810 18480
rect 4900 18240 5140 18480
rect 5230 18240 5470 18480
rect 5560 18240 5800 18480
rect 5890 18240 6130 18480
rect 6220 18240 6460 18480
rect 6550 18240 6790 18480
rect 6880 18240 7120 18480
rect -4670 17910 -4430 18150
rect -4340 17910 -4100 18150
rect -4010 17910 -3770 18150
rect -3680 17910 -3440 18150
rect -3350 17910 -3110 18150
rect -3020 17910 -2780 18150
rect -2690 17910 -2450 18150
rect -2360 17910 -2120 18150
rect -2030 17910 -1790 18150
rect -1700 17910 -1460 18150
rect -1370 17910 -1130 18150
rect -1040 17910 -800 18150
rect -710 17910 -470 18150
rect -380 17910 -140 18150
rect -50 17910 190 18150
rect 280 17910 520 18150
rect 610 17910 850 18150
rect 940 17910 1180 18150
rect 1270 17910 1510 18150
rect 1600 17910 1840 18150
rect 1930 17910 2170 18150
rect 2260 17910 2500 18150
rect 2590 17910 2830 18150
rect 2920 17910 3160 18150
rect 3250 17910 3490 18150
rect 3580 17910 3820 18150
rect 3910 17910 4150 18150
rect 4240 17910 4480 18150
rect 4570 17910 4810 18150
rect 4900 17910 5140 18150
rect 5230 17910 5470 18150
rect 5560 17910 5800 18150
rect 5890 17910 6130 18150
rect 6220 17910 6460 18150
rect 6550 17910 6790 18150
rect 6880 17910 7120 18150
rect -4670 17580 -4430 17820
rect -4340 17580 -4100 17820
rect -4010 17580 -3770 17820
rect -3680 17580 -3440 17820
rect -3350 17580 -3110 17820
rect -3020 17580 -2780 17820
rect -2690 17580 -2450 17820
rect -2360 17580 -2120 17820
rect -2030 17580 -1790 17820
rect -1700 17580 -1460 17820
rect -1370 17580 -1130 17820
rect -1040 17580 -800 17820
rect -710 17580 -470 17820
rect -380 17580 -140 17820
rect -50 17580 190 17820
rect 280 17580 520 17820
rect 610 17580 850 17820
rect 940 17580 1180 17820
rect 1270 17580 1510 17820
rect 1600 17580 1840 17820
rect 1930 17580 2170 17820
rect 2260 17580 2500 17820
rect 2590 17580 2830 17820
rect 2920 17580 3160 17820
rect 3250 17580 3490 17820
rect 3580 17580 3820 17820
rect 3910 17580 4150 17820
rect 4240 17580 4480 17820
rect 4570 17580 4810 17820
rect 4900 17580 5140 17820
rect 5230 17580 5470 17820
rect 5560 17580 5800 17820
rect 5890 17580 6130 17820
rect 6220 17580 6460 17820
rect 6550 17580 6790 17820
rect 6880 17580 7120 17820
rect -4670 17250 -4430 17490
rect -4340 17250 -4100 17490
rect -4010 17250 -3770 17490
rect -3680 17250 -3440 17490
rect -3350 17250 -3110 17490
rect -3020 17250 -2780 17490
rect -2690 17250 -2450 17490
rect -2360 17250 -2120 17490
rect -2030 17250 -1790 17490
rect -1700 17250 -1460 17490
rect -1370 17250 -1130 17490
rect -1040 17250 -800 17490
rect -710 17250 -470 17490
rect -380 17250 -140 17490
rect -50 17250 190 17490
rect 280 17250 520 17490
rect 610 17250 850 17490
rect 940 17250 1180 17490
rect 1270 17250 1510 17490
rect 1600 17250 1840 17490
rect 1930 17250 2170 17490
rect 2260 17250 2500 17490
rect 2590 17250 2830 17490
rect 2920 17250 3160 17490
rect 3250 17250 3490 17490
rect 3580 17250 3820 17490
rect 3910 17250 4150 17490
rect 4240 17250 4480 17490
rect 4570 17250 4810 17490
rect 4900 17250 5140 17490
rect 5230 17250 5470 17490
rect 5560 17250 5800 17490
rect 5890 17250 6130 17490
rect 6220 17250 6460 17490
rect 6550 17250 6790 17490
rect 6880 17250 7120 17490
rect -4670 16920 -4430 17160
rect -4340 16920 -4100 17160
rect -4010 16920 -3770 17160
rect -3680 16920 -3440 17160
rect -3350 16920 -3110 17160
rect -3020 16920 -2780 17160
rect -2690 16920 -2450 17160
rect -2360 16920 -2120 17160
rect -2030 16920 -1790 17160
rect -1700 16920 -1460 17160
rect -1370 16920 -1130 17160
rect -1040 16920 -800 17160
rect -710 16920 -470 17160
rect -380 16920 -140 17160
rect -50 16920 190 17160
rect 280 16920 520 17160
rect 610 16920 850 17160
rect 940 16920 1180 17160
rect 1270 16920 1510 17160
rect 1600 16920 1840 17160
rect 1930 16920 2170 17160
rect 2260 16920 2500 17160
rect 2590 16920 2830 17160
rect 2920 16920 3160 17160
rect 3250 16920 3490 17160
rect 3580 16920 3820 17160
rect 3910 16920 4150 17160
rect 4240 16920 4480 17160
rect 4570 16920 4810 17160
rect 4900 16920 5140 17160
rect 5230 16920 5470 17160
rect 5560 16920 5800 17160
rect 5890 16920 6130 17160
rect 6220 16920 6460 17160
rect 6550 16920 6790 17160
rect 6880 16920 7120 17160
rect -4670 16590 -4430 16830
rect -4340 16590 -4100 16830
rect -4010 16590 -3770 16830
rect -3680 16590 -3440 16830
rect -3350 16590 -3110 16830
rect -3020 16590 -2780 16830
rect -2690 16590 -2450 16830
rect -2360 16590 -2120 16830
rect -2030 16590 -1790 16830
rect -1700 16590 -1460 16830
rect -1370 16590 -1130 16830
rect -1040 16590 -800 16830
rect -710 16590 -470 16830
rect -380 16590 -140 16830
rect -50 16590 190 16830
rect 280 16590 520 16830
rect 610 16590 850 16830
rect 940 16590 1180 16830
rect 1270 16590 1510 16830
rect 1600 16590 1840 16830
rect 1930 16590 2170 16830
rect 2260 16590 2500 16830
rect 2590 16590 2830 16830
rect 2920 16590 3160 16830
rect 3250 16590 3490 16830
rect 3580 16590 3820 16830
rect 3910 16590 4150 16830
rect 4240 16590 4480 16830
rect 4570 16590 4810 16830
rect 4900 16590 5140 16830
rect 5230 16590 5470 16830
rect 5560 16590 5800 16830
rect 5890 16590 6130 16830
rect 6220 16590 6460 16830
rect 6550 16590 6790 16830
rect 6880 16590 7120 16830
rect -4670 16260 -4430 16500
rect -4340 16260 -4100 16500
rect -4010 16260 -3770 16500
rect -3680 16260 -3440 16500
rect -3350 16260 -3110 16500
rect -3020 16260 -2780 16500
rect -2690 16260 -2450 16500
rect -2360 16260 -2120 16500
rect -2030 16260 -1790 16500
rect -1700 16260 -1460 16500
rect -1370 16260 -1130 16500
rect -1040 16260 -800 16500
rect -710 16260 -470 16500
rect -380 16260 -140 16500
rect -50 16260 190 16500
rect 280 16260 520 16500
rect 610 16260 850 16500
rect 940 16260 1180 16500
rect 1270 16260 1510 16500
rect 1600 16260 1840 16500
rect 1930 16260 2170 16500
rect 2260 16260 2500 16500
rect 2590 16260 2830 16500
rect 2920 16260 3160 16500
rect 3250 16260 3490 16500
rect 3580 16260 3820 16500
rect 3910 16260 4150 16500
rect 4240 16260 4480 16500
rect 4570 16260 4810 16500
rect 4900 16260 5140 16500
rect 5230 16260 5470 16500
rect 5560 16260 5800 16500
rect 5890 16260 6130 16500
rect 6220 16260 6460 16500
rect 6550 16260 6790 16500
rect 6880 16260 7120 16500
rect -4670 15930 -4430 16170
rect -4340 15930 -4100 16170
rect -4010 15930 -3770 16170
rect -3680 15930 -3440 16170
rect -3350 15930 -3110 16170
rect -3020 15930 -2780 16170
rect -2690 15930 -2450 16170
rect -2360 15930 -2120 16170
rect -2030 15930 -1790 16170
rect -1700 15930 -1460 16170
rect -1370 15930 -1130 16170
rect -1040 15930 -800 16170
rect -710 15930 -470 16170
rect -380 15930 -140 16170
rect -50 15930 190 16170
rect 280 15930 520 16170
rect 610 15930 850 16170
rect 940 15930 1180 16170
rect 1270 15930 1510 16170
rect 1600 15930 1840 16170
rect 1930 15930 2170 16170
rect 2260 15930 2500 16170
rect 2590 15930 2830 16170
rect 2920 15930 3160 16170
rect 3250 15930 3490 16170
rect 3580 15930 3820 16170
rect 3910 15930 4150 16170
rect 4240 15930 4480 16170
rect 4570 15930 4810 16170
rect 4900 15930 5140 16170
rect 5230 15930 5470 16170
rect 5560 15930 5800 16170
rect 5890 15930 6130 16170
rect 6220 15930 6460 16170
rect 6550 15930 6790 16170
rect 6880 15930 7120 16170
rect -4670 15600 -4430 15840
rect -4340 15600 -4100 15840
rect -4010 15600 -3770 15840
rect -3680 15600 -3440 15840
rect -3350 15600 -3110 15840
rect -3020 15600 -2780 15840
rect -2690 15600 -2450 15840
rect -2360 15600 -2120 15840
rect -2030 15600 -1790 15840
rect -1700 15600 -1460 15840
rect -1370 15600 -1130 15840
rect -1040 15600 -800 15840
rect -710 15600 -470 15840
rect -380 15600 -140 15840
rect -50 15600 190 15840
rect 280 15600 520 15840
rect 610 15600 850 15840
rect 940 15600 1180 15840
rect 1270 15600 1510 15840
rect 1600 15600 1840 15840
rect 1930 15600 2170 15840
rect 2260 15600 2500 15840
rect 2590 15600 2830 15840
rect 2920 15600 3160 15840
rect 3250 15600 3490 15840
rect 3580 15600 3820 15840
rect 3910 15600 4150 15840
rect 4240 15600 4480 15840
rect 4570 15600 4810 15840
rect 4900 15600 5140 15840
rect 5230 15600 5470 15840
rect 5560 15600 5800 15840
rect 5890 15600 6130 15840
rect 6220 15600 6460 15840
rect 6550 15600 6790 15840
rect 6880 15600 7120 15840
rect -4670 15270 -4430 15510
rect -4340 15270 -4100 15510
rect -4010 15270 -3770 15510
rect -3680 15270 -3440 15510
rect -3350 15270 -3110 15510
rect -3020 15270 -2780 15510
rect -2690 15270 -2450 15510
rect -2360 15270 -2120 15510
rect -2030 15270 -1790 15510
rect -1700 15270 -1460 15510
rect -1370 15270 -1130 15510
rect -1040 15270 -800 15510
rect -710 15270 -470 15510
rect -380 15270 -140 15510
rect -50 15270 190 15510
rect 280 15270 520 15510
rect 610 15270 850 15510
rect 940 15270 1180 15510
rect 1270 15270 1510 15510
rect 1600 15270 1840 15510
rect 1930 15270 2170 15510
rect 2260 15270 2500 15510
rect 2590 15270 2830 15510
rect 2920 15270 3160 15510
rect 3250 15270 3490 15510
rect 3580 15270 3820 15510
rect 3910 15270 4150 15510
rect 4240 15270 4480 15510
rect 4570 15270 4810 15510
rect 4900 15270 5140 15510
rect 5230 15270 5470 15510
rect 5560 15270 5800 15510
rect 5890 15270 6130 15510
rect 6220 15270 6460 15510
rect 6550 15270 6790 15510
rect 6880 15270 7120 15510
rect -4670 14940 -4430 15180
rect -4340 14940 -4100 15180
rect -4010 14940 -3770 15180
rect -3680 14940 -3440 15180
rect -3350 14940 -3110 15180
rect -3020 14940 -2780 15180
rect -2690 14940 -2450 15180
rect -2360 14940 -2120 15180
rect -2030 14940 -1790 15180
rect -1700 14940 -1460 15180
rect -1370 14940 -1130 15180
rect -1040 14940 -800 15180
rect -710 14940 -470 15180
rect -380 14940 -140 15180
rect -50 14940 190 15180
rect 280 14940 520 15180
rect 610 14940 850 15180
rect 940 14940 1180 15180
rect 1270 14940 1510 15180
rect 1600 14940 1840 15180
rect 1930 14940 2170 15180
rect 2260 14940 2500 15180
rect 2590 14940 2830 15180
rect 2920 14940 3160 15180
rect 3250 14940 3490 15180
rect 3580 14940 3820 15180
rect 3910 14940 4150 15180
rect 4240 14940 4480 15180
rect 4570 14940 4810 15180
rect 4900 14940 5140 15180
rect 5230 14940 5470 15180
rect 5560 14940 5800 15180
rect 5890 14940 6130 15180
rect 6220 14940 6460 15180
rect 6550 14940 6790 15180
rect 6880 14940 7120 15180
rect -4670 14610 -4430 14850
rect -4340 14610 -4100 14850
rect -4010 14610 -3770 14850
rect -3680 14610 -3440 14850
rect -3350 14610 -3110 14850
rect -3020 14610 -2780 14850
rect -2690 14610 -2450 14850
rect -2360 14610 -2120 14850
rect -2030 14610 -1790 14850
rect -1700 14610 -1460 14850
rect -1370 14610 -1130 14850
rect -1040 14610 -800 14850
rect -710 14610 -470 14850
rect -380 14610 -140 14850
rect -50 14610 190 14850
rect 280 14610 520 14850
rect 610 14610 850 14850
rect 940 14610 1180 14850
rect 1270 14610 1510 14850
rect 1600 14610 1840 14850
rect 1930 14610 2170 14850
rect 2260 14610 2500 14850
rect 2590 14610 2830 14850
rect 2920 14610 3160 14850
rect 3250 14610 3490 14850
rect 3580 14610 3820 14850
rect 3910 14610 4150 14850
rect 4240 14610 4480 14850
rect 4570 14610 4810 14850
rect 4900 14610 5140 14850
rect 5230 14610 5470 14850
rect 5560 14610 5800 14850
rect 5890 14610 6130 14850
rect 6220 14610 6460 14850
rect 6550 14610 6790 14850
rect 6880 14610 7120 14850
rect -4670 14280 -4430 14520
rect -4340 14280 -4100 14520
rect -4010 14280 -3770 14520
rect -3680 14280 -3440 14520
rect -3350 14280 -3110 14520
rect -3020 14280 -2780 14520
rect -2690 14280 -2450 14520
rect -2360 14280 -2120 14520
rect -2030 14280 -1790 14520
rect -1700 14280 -1460 14520
rect -1370 14280 -1130 14520
rect -1040 14280 -800 14520
rect -710 14280 -470 14520
rect -380 14280 -140 14520
rect -50 14280 190 14520
rect 280 14280 520 14520
rect 610 14280 850 14520
rect 940 14280 1180 14520
rect 1270 14280 1510 14520
rect 1600 14280 1840 14520
rect 1930 14280 2170 14520
rect 2260 14280 2500 14520
rect 2590 14280 2830 14520
rect 2920 14280 3160 14520
rect 3250 14280 3490 14520
rect 3580 14280 3820 14520
rect 3910 14280 4150 14520
rect 4240 14280 4480 14520
rect 4570 14280 4810 14520
rect 4900 14280 5140 14520
rect 5230 14280 5470 14520
rect 5560 14280 5800 14520
rect 5890 14280 6130 14520
rect 6220 14280 6460 14520
rect 6550 14280 6790 14520
rect 6880 14280 7120 14520
rect -4670 13950 -4430 14190
rect -4340 13950 -4100 14190
rect -4010 13950 -3770 14190
rect -3680 13950 -3440 14190
rect -3350 13950 -3110 14190
rect -3020 13950 -2780 14190
rect -2690 13950 -2450 14190
rect -2360 13950 -2120 14190
rect -2030 13950 -1790 14190
rect -1700 13950 -1460 14190
rect -1370 13950 -1130 14190
rect -1040 13950 -800 14190
rect -710 13950 -470 14190
rect -380 13950 -140 14190
rect -50 13950 190 14190
rect 280 13950 520 14190
rect 610 13950 850 14190
rect 940 13950 1180 14190
rect 1270 13950 1510 14190
rect 1600 13950 1840 14190
rect 1930 13950 2170 14190
rect 2260 13950 2500 14190
rect 2590 13950 2830 14190
rect 2920 13950 3160 14190
rect 3250 13950 3490 14190
rect 3580 13950 3820 14190
rect 3910 13950 4150 14190
rect 4240 13950 4480 14190
rect 4570 13950 4810 14190
rect 4900 13950 5140 14190
rect 5230 13950 5470 14190
rect 5560 13950 5800 14190
rect 5890 13950 6130 14190
rect 6220 13950 6460 14190
rect 6550 13950 6790 14190
rect 6880 13950 7120 14190
rect -4670 13620 -4430 13860
rect -4340 13620 -4100 13860
rect -4010 13620 -3770 13860
rect -3680 13620 -3440 13860
rect -3350 13620 -3110 13860
rect -3020 13620 -2780 13860
rect -2690 13620 -2450 13860
rect -2360 13620 -2120 13860
rect -2030 13620 -1790 13860
rect -1700 13620 -1460 13860
rect -1370 13620 -1130 13860
rect -1040 13620 -800 13860
rect -710 13620 -470 13860
rect -380 13620 -140 13860
rect -50 13620 190 13860
rect 280 13620 520 13860
rect 610 13620 850 13860
rect 940 13620 1180 13860
rect 1270 13620 1510 13860
rect 1600 13620 1840 13860
rect 1930 13620 2170 13860
rect 2260 13620 2500 13860
rect 2590 13620 2830 13860
rect 2920 13620 3160 13860
rect 3250 13620 3490 13860
rect 3580 13620 3820 13860
rect 3910 13620 4150 13860
rect 4240 13620 4480 13860
rect 4570 13620 4810 13860
rect 4900 13620 5140 13860
rect 5230 13620 5470 13860
rect 5560 13620 5800 13860
rect 5890 13620 6130 13860
rect 6220 13620 6460 13860
rect 6550 13620 6790 13860
rect 6880 13620 7120 13860
rect -4670 13290 -4430 13530
rect -4340 13290 -4100 13530
rect -4010 13290 -3770 13530
rect -3680 13290 -3440 13530
rect -3350 13290 -3110 13530
rect -3020 13290 -2780 13530
rect -2690 13290 -2450 13530
rect -2360 13290 -2120 13530
rect -2030 13290 -1790 13530
rect -1700 13290 -1460 13530
rect -1370 13290 -1130 13530
rect -1040 13290 -800 13530
rect -710 13290 -470 13530
rect -380 13290 -140 13530
rect -50 13290 190 13530
rect 280 13290 520 13530
rect 610 13290 850 13530
rect 940 13290 1180 13530
rect 1270 13290 1510 13530
rect 1600 13290 1840 13530
rect 1930 13290 2170 13530
rect 2260 13290 2500 13530
rect 2590 13290 2830 13530
rect 2920 13290 3160 13530
rect 3250 13290 3490 13530
rect 3580 13290 3820 13530
rect 3910 13290 4150 13530
rect 4240 13290 4480 13530
rect 4570 13290 4810 13530
rect 4900 13290 5140 13530
rect 5230 13290 5470 13530
rect 5560 13290 5800 13530
rect 5890 13290 6130 13530
rect 6220 13290 6460 13530
rect 6550 13290 6790 13530
rect 6880 13290 7120 13530
rect -4670 12960 -4430 13200
rect -4340 12960 -4100 13200
rect -4010 12960 -3770 13200
rect -3680 12960 -3440 13200
rect -3350 12960 -3110 13200
rect -3020 12960 -2780 13200
rect -2690 12960 -2450 13200
rect -2360 12960 -2120 13200
rect -2030 12960 -1790 13200
rect -1700 12960 -1460 13200
rect -1370 12960 -1130 13200
rect -1040 12960 -800 13200
rect -710 12960 -470 13200
rect -380 12960 -140 13200
rect -50 12960 190 13200
rect 280 12960 520 13200
rect 610 12960 850 13200
rect 940 12960 1180 13200
rect 1270 12960 1510 13200
rect 1600 12960 1840 13200
rect 1930 12960 2170 13200
rect 2260 12960 2500 13200
rect 2590 12960 2830 13200
rect 2920 12960 3160 13200
rect 3250 12960 3490 13200
rect 3580 12960 3820 13200
rect 3910 12960 4150 13200
rect 4240 12960 4480 13200
rect 4570 12960 4810 13200
rect 4900 12960 5140 13200
rect 5230 12960 5470 13200
rect 5560 12960 5800 13200
rect 5890 12960 6130 13200
rect 6220 12960 6460 13200
rect 6550 12960 6790 13200
rect 6880 12960 7120 13200
rect -4670 12630 -4430 12870
rect -4340 12630 -4100 12870
rect -4010 12630 -3770 12870
rect -3680 12630 -3440 12870
rect -3350 12630 -3110 12870
rect -3020 12630 -2780 12870
rect -2690 12630 -2450 12870
rect -2360 12630 -2120 12870
rect -2030 12630 -1790 12870
rect -1700 12630 -1460 12870
rect -1370 12630 -1130 12870
rect -1040 12630 -800 12870
rect -710 12630 -470 12870
rect -380 12630 -140 12870
rect -50 12630 190 12870
rect 280 12630 520 12870
rect 610 12630 850 12870
rect 940 12630 1180 12870
rect 1270 12630 1510 12870
rect 1600 12630 1840 12870
rect 1930 12630 2170 12870
rect 2260 12630 2500 12870
rect 2590 12630 2830 12870
rect 2920 12630 3160 12870
rect 3250 12630 3490 12870
rect 3580 12630 3820 12870
rect 3910 12630 4150 12870
rect 4240 12630 4480 12870
rect 4570 12630 4810 12870
rect 4900 12630 5140 12870
rect 5230 12630 5470 12870
rect 5560 12630 5800 12870
rect 5890 12630 6130 12870
rect 6220 12630 6460 12870
rect 6550 12630 6790 12870
rect 6880 12630 7120 12870
rect -4670 12300 -4430 12540
rect -4340 12300 -4100 12540
rect -4010 12300 -3770 12540
rect -3680 12300 -3440 12540
rect -3350 12300 -3110 12540
rect -3020 12300 -2780 12540
rect -2690 12300 -2450 12540
rect -2360 12300 -2120 12540
rect -2030 12300 -1790 12540
rect -1700 12300 -1460 12540
rect -1370 12300 -1130 12540
rect -1040 12300 -800 12540
rect -710 12300 -470 12540
rect -380 12300 -140 12540
rect -50 12300 190 12540
rect 280 12300 520 12540
rect 610 12300 850 12540
rect 940 12300 1180 12540
rect 1270 12300 1510 12540
rect 1600 12300 1840 12540
rect 1930 12300 2170 12540
rect 2260 12300 2500 12540
rect 2590 12300 2830 12540
rect 2920 12300 3160 12540
rect 3250 12300 3490 12540
rect 3580 12300 3820 12540
rect 3910 12300 4150 12540
rect 4240 12300 4480 12540
rect 4570 12300 4810 12540
rect 4900 12300 5140 12540
rect 5230 12300 5470 12540
rect 5560 12300 5800 12540
rect 5890 12300 6130 12540
rect 6220 12300 6460 12540
rect 6550 12300 6790 12540
rect 6880 12300 7120 12540
rect -4670 11970 -4430 12210
rect -4340 11970 -4100 12210
rect -4010 11970 -3770 12210
rect -3680 11970 -3440 12210
rect -3350 11970 -3110 12210
rect -3020 11970 -2780 12210
rect -2690 11970 -2450 12210
rect -2360 11970 -2120 12210
rect -2030 11970 -1790 12210
rect -1700 11970 -1460 12210
rect -1370 11970 -1130 12210
rect -1040 11970 -800 12210
rect -710 11970 -470 12210
rect -380 11970 -140 12210
rect -50 11970 190 12210
rect 280 11970 520 12210
rect 610 11970 850 12210
rect 940 11970 1180 12210
rect 1270 11970 1510 12210
rect 1600 11970 1840 12210
rect 1930 11970 2170 12210
rect 2260 11970 2500 12210
rect 2590 11970 2830 12210
rect 2920 11970 3160 12210
rect 3250 11970 3490 12210
rect 3580 11970 3820 12210
rect 3910 11970 4150 12210
rect 4240 11970 4480 12210
rect 4570 11970 4810 12210
rect 4900 11970 5140 12210
rect 5230 11970 5470 12210
rect 5560 11970 5800 12210
rect 5890 11970 6130 12210
rect 6220 11970 6460 12210
rect 6550 11970 6790 12210
rect 6880 11970 7120 12210
rect -4670 11640 -4430 11880
rect -4340 11640 -4100 11880
rect -4010 11640 -3770 11880
rect -3680 11640 -3440 11880
rect -3350 11640 -3110 11880
rect -3020 11640 -2780 11880
rect -2690 11640 -2450 11880
rect -2360 11640 -2120 11880
rect -2030 11640 -1790 11880
rect -1700 11640 -1460 11880
rect -1370 11640 -1130 11880
rect -1040 11640 -800 11880
rect -710 11640 -470 11880
rect -380 11640 -140 11880
rect -50 11640 190 11880
rect 280 11640 520 11880
rect 610 11640 850 11880
rect 940 11640 1180 11880
rect 1270 11640 1510 11880
rect 1600 11640 1840 11880
rect 1930 11640 2170 11880
rect 2260 11640 2500 11880
rect 2590 11640 2830 11880
rect 2920 11640 3160 11880
rect 3250 11640 3490 11880
rect 3580 11640 3820 11880
rect 3910 11640 4150 11880
rect 4240 11640 4480 11880
rect 4570 11640 4810 11880
rect 4900 11640 5140 11880
rect 5230 11640 5470 11880
rect 5560 11640 5800 11880
rect 5890 11640 6130 11880
rect 6220 11640 6460 11880
rect 6550 11640 6790 11880
rect 6880 11640 7120 11880
rect -4670 11310 -4430 11550
rect -4340 11310 -4100 11550
rect -4010 11310 -3770 11550
rect -3680 11310 -3440 11550
rect -3350 11310 -3110 11550
rect -3020 11310 -2780 11550
rect -2690 11310 -2450 11550
rect -2360 11310 -2120 11550
rect -2030 11310 -1790 11550
rect -1700 11310 -1460 11550
rect -1370 11310 -1130 11550
rect -1040 11310 -800 11550
rect -710 11310 -470 11550
rect -380 11310 -140 11550
rect -50 11310 190 11550
rect 280 11310 520 11550
rect 610 11310 850 11550
rect 940 11310 1180 11550
rect 1270 11310 1510 11550
rect 1600 11310 1840 11550
rect 1930 11310 2170 11550
rect 2260 11310 2500 11550
rect 2590 11310 2830 11550
rect 2920 11310 3160 11550
rect 3250 11310 3490 11550
rect 3580 11310 3820 11550
rect 3910 11310 4150 11550
rect 4240 11310 4480 11550
rect 4570 11310 4810 11550
rect 4900 11310 5140 11550
rect 5230 11310 5470 11550
rect 5560 11310 5800 11550
rect 5890 11310 6130 11550
rect 6220 11310 6460 11550
rect 6550 11310 6790 11550
rect 6880 11310 7120 11550
rect -4670 10980 -4430 11220
rect -4340 10980 -4100 11220
rect -4010 10980 -3770 11220
rect -3680 10980 -3440 11220
rect -3350 10980 -3110 11220
rect -3020 10980 -2780 11220
rect -2690 10980 -2450 11220
rect -2360 10980 -2120 11220
rect -2030 10980 -1790 11220
rect -1700 10980 -1460 11220
rect -1370 10980 -1130 11220
rect -1040 10980 -800 11220
rect -710 10980 -470 11220
rect -380 10980 -140 11220
rect -50 10980 190 11220
rect 280 10980 520 11220
rect 610 10980 850 11220
rect 940 10980 1180 11220
rect 1270 10980 1510 11220
rect 1600 10980 1840 11220
rect 1930 10980 2170 11220
rect 2260 10980 2500 11220
rect 2590 10980 2830 11220
rect 2920 10980 3160 11220
rect 3250 10980 3490 11220
rect 3580 10980 3820 11220
rect 3910 10980 4150 11220
rect 4240 10980 4480 11220
rect 4570 10980 4810 11220
rect 4900 10980 5140 11220
rect 5230 10980 5470 11220
rect 5560 10980 5800 11220
rect 5890 10980 6130 11220
rect 6220 10980 6460 11220
rect 6550 10980 6790 11220
rect 6880 10980 7120 11220
rect -4670 10650 -4430 10890
rect -4340 10650 -4100 10890
rect -4010 10650 -3770 10890
rect -3680 10650 -3440 10890
rect -3350 10650 -3110 10890
rect -3020 10650 -2780 10890
rect -2690 10650 -2450 10890
rect -2360 10650 -2120 10890
rect -2030 10650 -1790 10890
rect -1700 10650 -1460 10890
rect -1370 10650 -1130 10890
rect -1040 10650 -800 10890
rect -710 10650 -470 10890
rect -380 10650 -140 10890
rect -50 10650 190 10890
rect 280 10650 520 10890
rect 610 10650 850 10890
rect 940 10650 1180 10890
rect 1270 10650 1510 10890
rect 1600 10650 1840 10890
rect 1930 10650 2170 10890
rect 2260 10650 2500 10890
rect 2590 10650 2830 10890
rect 2920 10650 3160 10890
rect 3250 10650 3490 10890
rect 3580 10650 3820 10890
rect 3910 10650 4150 10890
rect 4240 10650 4480 10890
rect 4570 10650 4810 10890
rect 4900 10650 5140 10890
rect 5230 10650 5470 10890
rect 5560 10650 5800 10890
rect 5890 10650 6130 10890
rect 6220 10650 6460 10890
rect 6550 10650 6790 10890
rect 6880 10650 7120 10890
rect -4670 10320 -4430 10560
rect -4340 10320 -4100 10560
rect -4010 10320 -3770 10560
rect -3680 10320 -3440 10560
rect -3350 10320 -3110 10560
rect -3020 10320 -2780 10560
rect -2690 10320 -2450 10560
rect -2360 10320 -2120 10560
rect -2030 10320 -1790 10560
rect -1700 10320 -1460 10560
rect -1370 10320 -1130 10560
rect -1040 10320 -800 10560
rect -710 10320 -470 10560
rect -380 10320 -140 10560
rect -50 10320 190 10560
rect 280 10320 520 10560
rect 610 10320 850 10560
rect 940 10320 1180 10560
rect 1270 10320 1510 10560
rect 1600 10320 1840 10560
rect 1930 10320 2170 10560
rect 2260 10320 2500 10560
rect 2590 10320 2830 10560
rect 2920 10320 3160 10560
rect 3250 10320 3490 10560
rect 3580 10320 3820 10560
rect 3910 10320 4150 10560
rect 4240 10320 4480 10560
rect 4570 10320 4810 10560
rect 4900 10320 5140 10560
rect 5230 10320 5470 10560
rect 5560 10320 5800 10560
rect 5890 10320 6130 10560
rect 6220 10320 6460 10560
rect 6550 10320 6790 10560
rect 6880 10320 7120 10560
rect -4670 9990 -4430 10230
rect -4340 9990 -4100 10230
rect -4010 9990 -3770 10230
rect -3680 9990 -3440 10230
rect -3350 9990 -3110 10230
rect -3020 9990 -2780 10230
rect -2690 9990 -2450 10230
rect -2360 9990 -2120 10230
rect -2030 9990 -1790 10230
rect -1700 9990 -1460 10230
rect -1370 9990 -1130 10230
rect -1040 9990 -800 10230
rect -710 9990 -470 10230
rect -380 9990 -140 10230
rect -50 9990 190 10230
rect 280 9990 520 10230
rect 610 9990 850 10230
rect 940 9990 1180 10230
rect 1270 9990 1510 10230
rect 1600 9990 1840 10230
rect 1930 9990 2170 10230
rect 2260 9990 2500 10230
rect 2590 9990 2830 10230
rect 2920 9990 3160 10230
rect 3250 9990 3490 10230
rect 3580 9990 3820 10230
rect 3910 9990 4150 10230
rect 4240 9990 4480 10230
rect 4570 9990 4810 10230
rect 4900 9990 5140 10230
rect 5230 9990 5470 10230
rect 5560 9990 5800 10230
rect 5890 9990 6130 10230
rect 6220 9990 6460 10230
rect 6550 9990 6790 10230
rect 6880 9990 7120 10230
rect -4670 9660 -4430 9900
rect -4340 9660 -4100 9900
rect -4010 9660 -3770 9900
rect -3680 9660 -3440 9900
rect -3350 9660 -3110 9900
rect -3020 9660 -2780 9900
rect -2690 9660 -2450 9900
rect -2360 9660 -2120 9900
rect -2030 9660 -1790 9900
rect -1700 9660 -1460 9900
rect -1370 9660 -1130 9900
rect -1040 9660 -800 9900
rect -710 9660 -470 9900
rect -380 9660 -140 9900
rect -50 9660 190 9900
rect 280 9660 520 9900
rect 610 9660 850 9900
rect 940 9660 1180 9900
rect 1270 9660 1510 9900
rect 1600 9660 1840 9900
rect 1930 9660 2170 9900
rect 2260 9660 2500 9900
rect 2590 9660 2830 9900
rect 2920 9660 3160 9900
rect 3250 9660 3490 9900
rect 3580 9660 3820 9900
rect 3910 9660 4150 9900
rect 4240 9660 4480 9900
rect 4570 9660 4810 9900
rect 4900 9660 5140 9900
rect 5230 9660 5470 9900
rect 5560 9660 5800 9900
rect 5890 9660 6130 9900
rect 6220 9660 6460 9900
rect 6550 9660 6790 9900
rect 6880 9660 7120 9900
rect -4670 9330 -4430 9570
rect -4340 9330 -4100 9570
rect -4010 9330 -3770 9570
rect -3680 9330 -3440 9570
rect -3350 9330 -3110 9570
rect -3020 9330 -2780 9570
rect -2690 9330 -2450 9570
rect -2360 9330 -2120 9570
rect -2030 9330 -1790 9570
rect -1700 9330 -1460 9570
rect -1370 9330 -1130 9570
rect -1040 9330 -800 9570
rect -710 9330 -470 9570
rect -380 9330 -140 9570
rect -50 9330 190 9570
rect 280 9330 520 9570
rect 610 9330 850 9570
rect 940 9330 1180 9570
rect 1270 9330 1510 9570
rect 1600 9330 1840 9570
rect 1930 9330 2170 9570
rect 2260 9330 2500 9570
rect 2590 9330 2830 9570
rect 2920 9330 3160 9570
rect 3250 9330 3490 9570
rect 3580 9330 3820 9570
rect 3910 9330 4150 9570
rect 4240 9330 4480 9570
rect 4570 9330 4810 9570
rect 4900 9330 5140 9570
rect 5230 9330 5470 9570
rect 5560 9330 5800 9570
rect 5890 9330 6130 9570
rect 6220 9330 6460 9570
rect 6550 9330 6790 9570
rect 6880 9330 7120 9570
rect -4670 9000 -4430 9240
rect -4340 9000 -4100 9240
rect -4010 9000 -3770 9240
rect -3680 9000 -3440 9240
rect -3350 9000 -3110 9240
rect -3020 9000 -2780 9240
rect -2690 9000 -2450 9240
rect -2360 9000 -2120 9240
rect -2030 9000 -1790 9240
rect -1700 9000 -1460 9240
rect -1370 9000 -1130 9240
rect -1040 9000 -800 9240
rect -710 9000 -470 9240
rect -380 9000 -140 9240
rect -50 9000 190 9240
rect 280 9000 520 9240
rect 610 9000 850 9240
rect 940 9000 1180 9240
rect 1270 9000 1510 9240
rect 1600 9000 1840 9240
rect 1930 9000 2170 9240
rect 2260 9000 2500 9240
rect 2590 9000 2830 9240
rect 2920 9000 3160 9240
rect 3250 9000 3490 9240
rect 3580 9000 3820 9240
rect 3910 9000 4150 9240
rect 4240 9000 4480 9240
rect 4570 9000 4810 9240
rect 4900 9000 5140 9240
rect 5230 9000 5470 9240
rect 5560 9000 5800 9240
rect 5890 9000 6130 9240
rect 6220 9000 6460 9240
rect 6550 9000 6790 9240
rect 6880 9000 7120 9240
rect 7780 20550 8020 20790
rect 8110 20550 8350 20790
rect 8440 20550 8680 20790
rect 8770 20550 9010 20790
rect 9100 20550 9340 20790
rect 9430 20550 9670 20790
rect 9760 20550 10000 20790
rect 10090 20550 10330 20790
rect 10420 20550 10660 20790
rect 10750 20550 10990 20790
rect 11080 20550 11320 20790
rect 11410 20550 11650 20790
rect 11740 20550 11980 20790
rect 12070 20550 12310 20790
rect 12400 20550 12640 20790
rect 12730 20550 12970 20790
rect 13060 20550 13300 20790
rect 13390 20550 13630 20790
rect 13720 20550 13960 20790
rect 14050 20550 14290 20790
rect 14380 20550 14620 20790
rect 14710 20550 14950 20790
rect 15040 20550 15280 20790
rect 15370 20550 15610 20790
rect 15700 20550 15940 20790
rect 16030 20550 16270 20790
rect 16360 20550 16600 20790
rect 16690 20550 16930 20790
rect 17020 20550 17260 20790
rect 17350 20550 17590 20790
rect 17680 20550 17920 20790
rect 18010 20550 18250 20790
rect 18340 20550 18580 20790
rect 18670 20550 18910 20790
rect 19000 20550 19240 20790
rect 19330 20550 19570 20790
rect 7780 20220 8020 20460
rect 8110 20220 8350 20460
rect 8440 20220 8680 20460
rect 8770 20220 9010 20460
rect 9100 20220 9340 20460
rect 9430 20220 9670 20460
rect 9760 20220 10000 20460
rect 10090 20220 10330 20460
rect 10420 20220 10660 20460
rect 10750 20220 10990 20460
rect 11080 20220 11320 20460
rect 11410 20220 11650 20460
rect 11740 20220 11980 20460
rect 12070 20220 12310 20460
rect 12400 20220 12640 20460
rect 12730 20220 12970 20460
rect 13060 20220 13300 20460
rect 13390 20220 13630 20460
rect 13720 20220 13960 20460
rect 14050 20220 14290 20460
rect 14380 20220 14620 20460
rect 14710 20220 14950 20460
rect 15040 20220 15280 20460
rect 15370 20220 15610 20460
rect 15700 20220 15940 20460
rect 16030 20220 16270 20460
rect 16360 20220 16600 20460
rect 16690 20220 16930 20460
rect 17020 20220 17260 20460
rect 17350 20220 17590 20460
rect 17680 20220 17920 20460
rect 18010 20220 18250 20460
rect 18340 20220 18580 20460
rect 18670 20220 18910 20460
rect 19000 20220 19240 20460
rect 19330 20220 19570 20460
rect 7780 19890 8020 20130
rect 8110 19890 8350 20130
rect 8440 19890 8680 20130
rect 8770 19890 9010 20130
rect 9100 19890 9340 20130
rect 9430 19890 9670 20130
rect 9760 19890 10000 20130
rect 10090 19890 10330 20130
rect 10420 19890 10660 20130
rect 10750 19890 10990 20130
rect 11080 19890 11320 20130
rect 11410 19890 11650 20130
rect 11740 19890 11980 20130
rect 12070 19890 12310 20130
rect 12400 19890 12640 20130
rect 12730 19890 12970 20130
rect 13060 19890 13300 20130
rect 13390 19890 13630 20130
rect 13720 19890 13960 20130
rect 14050 19890 14290 20130
rect 14380 19890 14620 20130
rect 14710 19890 14950 20130
rect 15040 19890 15280 20130
rect 15370 19890 15610 20130
rect 15700 19890 15940 20130
rect 16030 19890 16270 20130
rect 16360 19890 16600 20130
rect 16690 19890 16930 20130
rect 17020 19890 17260 20130
rect 17350 19890 17590 20130
rect 17680 19890 17920 20130
rect 18010 19890 18250 20130
rect 18340 19890 18580 20130
rect 18670 19890 18910 20130
rect 19000 19890 19240 20130
rect 19330 19890 19570 20130
rect 7780 19560 8020 19800
rect 8110 19560 8350 19800
rect 8440 19560 8680 19800
rect 8770 19560 9010 19800
rect 9100 19560 9340 19800
rect 9430 19560 9670 19800
rect 9760 19560 10000 19800
rect 10090 19560 10330 19800
rect 10420 19560 10660 19800
rect 10750 19560 10990 19800
rect 11080 19560 11320 19800
rect 11410 19560 11650 19800
rect 11740 19560 11980 19800
rect 12070 19560 12310 19800
rect 12400 19560 12640 19800
rect 12730 19560 12970 19800
rect 13060 19560 13300 19800
rect 13390 19560 13630 19800
rect 13720 19560 13960 19800
rect 14050 19560 14290 19800
rect 14380 19560 14620 19800
rect 14710 19560 14950 19800
rect 15040 19560 15280 19800
rect 15370 19560 15610 19800
rect 15700 19560 15940 19800
rect 16030 19560 16270 19800
rect 16360 19560 16600 19800
rect 16690 19560 16930 19800
rect 17020 19560 17260 19800
rect 17350 19560 17590 19800
rect 17680 19560 17920 19800
rect 18010 19560 18250 19800
rect 18340 19560 18580 19800
rect 18670 19560 18910 19800
rect 19000 19560 19240 19800
rect 19330 19560 19570 19800
rect 7780 19230 8020 19470
rect 8110 19230 8350 19470
rect 8440 19230 8680 19470
rect 8770 19230 9010 19470
rect 9100 19230 9340 19470
rect 9430 19230 9670 19470
rect 9760 19230 10000 19470
rect 10090 19230 10330 19470
rect 10420 19230 10660 19470
rect 10750 19230 10990 19470
rect 11080 19230 11320 19470
rect 11410 19230 11650 19470
rect 11740 19230 11980 19470
rect 12070 19230 12310 19470
rect 12400 19230 12640 19470
rect 12730 19230 12970 19470
rect 13060 19230 13300 19470
rect 13390 19230 13630 19470
rect 13720 19230 13960 19470
rect 14050 19230 14290 19470
rect 14380 19230 14620 19470
rect 14710 19230 14950 19470
rect 15040 19230 15280 19470
rect 15370 19230 15610 19470
rect 15700 19230 15940 19470
rect 16030 19230 16270 19470
rect 16360 19230 16600 19470
rect 16690 19230 16930 19470
rect 17020 19230 17260 19470
rect 17350 19230 17590 19470
rect 17680 19230 17920 19470
rect 18010 19230 18250 19470
rect 18340 19230 18580 19470
rect 18670 19230 18910 19470
rect 19000 19230 19240 19470
rect 19330 19230 19570 19470
rect 7780 18900 8020 19140
rect 8110 18900 8350 19140
rect 8440 18900 8680 19140
rect 8770 18900 9010 19140
rect 9100 18900 9340 19140
rect 9430 18900 9670 19140
rect 9760 18900 10000 19140
rect 10090 18900 10330 19140
rect 10420 18900 10660 19140
rect 10750 18900 10990 19140
rect 11080 18900 11320 19140
rect 11410 18900 11650 19140
rect 11740 18900 11980 19140
rect 12070 18900 12310 19140
rect 12400 18900 12640 19140
rect 12730 18900 12970 19140
rect 13060 18900 13300 19140
rect 13390 18900 13630 19140
rect 13720 18900 13960 19140
rect 14050 18900 14290 19140
rect 14380 18900 14620 19140
rect 14710 18900 14950 19140
rect 15040 18900 15280 19140
rect 15370 18900 15610 19140
rect 15700 18900 15940 19140
rect 16030 18900 16270 19140
rect 16360 18900 16600 19140
rect 16690 18900 16930 19140
rect 17020 18900 17260 19140
rect 17350 18900 17590 19140
rect 17680 18900 17920 19140
rect 18010 18900 18250 19140
rect 18340 18900 18580 19140
rect 18670 18900 18910 19140
rect 19000 18900 19240 19140
rect 19330 18900 19570 19140
rect 7780 18570 8020 18810
rect 8110 18570 8350 18810
rect 8440 18570 8680 18810
rect 8770 18570 9010 18810
rect 9100 18570 9340 18810
rect 9430 18570 9670 18810
rect 9760 18570 10000 18810
rect 10090 18570 10330 18810
rect 10420 18570 10660 18810
rect 10750 18570 10990 18810
rect 11080 18570 11320 18810
rect 11410 18570 11650 18810
rect 11740 18570 11980 18810
rect 12070 18570 12310 18810
rect 12400 18570 12640 18810
rect 12730 18570 12970 18810
rect 13060 18570 13300 18810
rect 13390 18570 13630 18810
rect 13720 18570 13960 18810
rect 14050 18570 14290 18810
rect 14380 18570 14620 18810
rect 14710 18570 14950 18810
rect 15040 18570 15280 18810
rect 15370 18570 15610 18810
rect 15700 18570 15940 18810
rect 16030 18570 16270 18810
rect 16360 18570 16600 18810
rect 16690 18570 16930 18810
rect 17020 18570 17260 18810
rect 17350 18570 17590 18810
rect 17680 18570 17920 18810
rect 18010 18570 18250 18810
rect 18340 18570 18580 18810
rect 18670 18570 18910 18810
rect 19000 18570 19240 18810
rect 19330 18570 19570 18810
rect 7780 18240 8020 18480
rect 8110 18240 8350 18480
rect 8440 18240 8680 18480
rect 8770 18240 9010 18480
rect 9100 18240 9340 18480
rect 9430 18240 9670 18480
rect 9760 18240 10000 18480
rect 10090 18240 10330 18480
rect 10420 18240 10660 18480
rect 10750 18240 10990 18480
rect 11080 18240 11320 18480
rect 11410 18240 11650 18480
rect 11740 18240 11980 18480
rect 12070 18240 12310 18480
rect 12400 18240 12640 18480
rect 12730 18240 12970 18480
rect 13060 18240 13300 18480
rect 13390 18240 13630 18480
rect 13720 18240 13960 18480
rect 14050 18240 14290 18480
rect 14380 18240 14620 18480
rect 14710 18240 14950 18480
rect 15040 18240 15280 18480
rect 15370 18240 15610 18480
rect 15700 18240 15940 18480
rect 16030 18240 16270 18480
rect 16360 18240 16600 18480
rect 16690 18240 16930 18480
rect 17020 18240 17260 18480
rect 17350 18240 17590 18480
rect 17680 18240 17920 18480
rect 18010 18240 18250 18480
rect 18340 18240 18580 18480
rect 18670 18240 18910 18480
rect 19000 18240 19240 18480
rect 19330 18240 19570 18480
rect 7780 17910 8020 18150
rect 8110 17910 8350 18150
rect 8440 17910 8680 18150
rect 8770 17910 9010 18150
rect 9100 17910 9340 18150
rect 9430 17910 9670 18150
rect 9760 17910 10000 18150
rect 10090 17910 10330 18150
rect 10420 17910 10660 18150
rect 10750 17910 10990 18150
rect 11080 17910 11320 18150
rect 11410 17910 11650 18150
rect 11740 17910 11980 18150
rect 12070 17910 12310 18150
rect 12400 17910 12640 18150
rect 12730 17910 12970 18150
rect 13060 17910 13300 18150
rect 13390 17910 13630 18150
rect 13720 17910 13960 18150
rect 14050 17910 14290 18150
rect 14380 17910 14620 18150
rect 14710 17910 14950 18150
rect 15040 17910 15280 18150
rect 15370 17910 15610 18150
rect 15700 17910 15940 18150
rect 16030 17910 16270 18150
rect 16360 17910 16600 18150
rect 16690 17910 16930 18150
rect 17020 17910 17260 18150
rect 17350 17910 17590 18150
rect 17680 17910 17920 18150
rect 18010 17910 18250 18150
rect 18340 17910 18580 18150
rect 18670 17910 18910 18150
rect 19000 17910 19240 18150
rect 19330 17910 19570 18150
rect 7780 17580 8020 17820
rect 8110 17580 8350 17820
rect 8440 17580 8680 17820
rect 8770 17580 9010 17820
rect 9100 17580 9340 17820
rect 9430 17580 9670 17820
rect 9760 17580 10000 17820
rect 10090 17580 10330 17820
rect 10420 17580 10660 17820
rect 10750 17580 10990 17820
rect 11080 17580 11320 17820
rect 11410 17580 11650 17820
rect 11740 17580 11980 17820
rect 12070 17580 12310 17820
rect 12400 17580 12640 17820
rect 12730 17580 12970 17820
rect 13060 17580 13300 17820
rect 13390 17580 13630 17820
rect 13720 17580 13960 17820
rect 14050 17580 14290 17820
rect 14380 17580 14620 17820
rect 14710 17580 14950 17820
rect 15040 17580 15280 17820
rect 15370 17580 15610 17820
rect 15700 17580 15940 17820
rect 16030 17580 16270 17820
rect 16360 17580 16600 17820
rect 16690 17580 16930 17820
rect 17020 17580 17260 17820
rect 17350 17580 17590 17820
rect 17680 17580 17920 17820
rect 18010 17580 18250 17820
rect 18340 17580 18580 17820
rect 18670 17580 18910 17820
rect 19000 17580 19240 17820
rect 19330 17580 19570 17820
rect 7780 17250 8020 17490
rect 8110 17250 8350 17490
rect 8440 17250 8680 17490
rect 8770 17250 9010 17490
rect 9100 17250 9340 17490
rect 9430 17250 9670 17490
rect 9760 17250 10000 17490
rect 10090 17250 10330 17490
rect 10420 17250 10660 17490
rect 10750 17250 10990 17490
rect 11080 17250 11320 17490
rect 11410 17250 11650 17490
rect 11740 17250 11980 17490
rect 12070 17250 12310 17490
rect 12400 17250 12640 17490
rect 12730 17250 12970 17490
rect 13060 17250 13300 17490
rect 13390 17250 13630 17490
rect 13720 17250 13960 17490
rect 14050 17250 14290 17490
rect 14380 17250 14620 17490
rect 14710 17250 14950 17490
rect 15040 17250 15280 17490
rect 15370 17250 15610 17490
rect 15700 17250 15940 17490
rect 16030 17250 16270 17490
rect 16360 17250 16600 17490
rect 16690 17250 16930 17490
rect 17020 17250 17260 17490
rect 17350 17250 17590 17490
rect 17680 17250 17920 17490
rect 18010 17250 18250 17490
rect 18340 17250 18580 17490
rect 18670 17250 18910 17490
rect 19000 17250 19240 17490
rect 19330 17250 19570 17490
rect 7780 16920 8020 17160
rect 8110 16920 8350 17160
rect 8440 16920 8680 17160
rect 8770 16920 9010 17160
rect 9100 16920 9340 17160
rect 9430 16920 9670 17160
rect 9760 16920 10000 17160
rect 10090 16920 10330 17160
rect 10420 16920 10660 17160
rect 10750 16920 10990 17160
rect 11080 16920 11320 17160
rect 11410 16920 11650 17160
rect 11740 16920 11980 17160
rect 12070 16920 12310 17160
rect 12400 16920 12640 17160
rect 12730 16920 12970 17160
rect 13060 16920 13300 17160
rect 13390 16920 13630 17160
rect 13720 16920 13960 17160
rect 14050 16920 14290 17160
rect 14380 16920 14620 17160
rect 14710 16920 14950 17160
rect 15040 16920 15280 17160
rect 15370 16920 15610 17160
rect 15700 16920 15940 17160
rect 16030 16920 16270 17160
rect 16360 16920 16600 17160
rect 16690 16920 16930 17160
rect 17020 16920 17260 17160
rect 17350 16920 17590 17160
rect 17680 16920 17920 17160
rect 18010 16920 18250 17160
rect 18340 16920 18580 17160
rect 18670 16920 18910 17160
rect 19000 16920 19240 17160
rect 19330 16920 19570 17160
rect 7780 16590 8020 16830
rect 8110 16590 8350 16830
rect 8440 16590 8680 16830
rect 8770 16590 9010 16830
rect 9100 16590 9340 16830
rect 9430 16590 9670 16830
rect 9760 16590 10000 16830
rect 10090 16590 10330 16830
rect 10420 16590 10660 16830
rect 10750 16590 10990 16830
rect 11080 16590 11320 16830
rect 11410 16590 11650 16830
rect 11740 16590 11980 16830
rect 12070 16590 12310 16830
rect 12400 16590 12640 16830
rect 12730 16590 12970 16830
rect 13060 16590 13300 16830
rect 13390 16590 13630 16830
rect 13720 16590 13960 16830
rect 14050 16590 14290 16830
rect 14380 16590 14620 16830
rect 14710 16590 14950 16830
rect 15040 16590 15280 16830
rect 15370 16590 15610 16830
rect 15700 16590 15940 16830
rect 16030 16590 16270 16830
rect 16360 16590 16600 16830
rect 16690 16590 16930 16830
rect 17020 16590 17260 16830
rect 17350 16590 17590 16830
rect 17680 16590 17920 16830
rect 18010 16590 18250 16830
rect 18340 16590 18580 16830
rect 18670 16590 18910 16830
rect 19000 16590 19240 16830
rect 19330 16590 19570 16830
rect 7780 16260 8020 16500
rect 8110 16260 8350 16500
rect 8440 16260 8680 16500
rect 8770 16260 9010 16500
rect 9100 16260 9340 16500
rect 9430 16260 9670 16500
rect 9760 16260 10000 16500
rect 10090 16260 10330 16500
rect 10420 16260 10660 16500
rect 10750 16260 10990 16500
rect 11080 16260 11320 16500
rect 11410 16260 11650 16500
rect 11740 16260 11980 16500
rect 12070 16260 12310 16500
rect 12400 16260 12640 16500
rect 12730 16260 12970 16500
rect 13060 16260 13300 16500
rect 13390 16260 13630 16500
rect 13720 16260 13960 16500
rect 14050 16260 14290 16500
rect 14380 16260 14620 16500
rect 14710 16260 14950 16500
rect 15040 16260 15280 16500
rect 15370 16260 15610 16500
rect 15700 16260 15940 16500
rect 16030 16260 16270 16500
rect 16360 16260 16600 16500
rect 16690 16260 16930 16500
rect 17020 16260 17260 16500
rect 17350 16260 17590 16500
rect 17680 16260 17920 16500
rect 18010 16260 18250 16500
rect 18340 16260 18580 16500
rect 18670 16260 18910 16500
rect 19000 16260 19240 16500
rect 19330 16260 19570 16500
rect 7780 15930 8020 16170
rect 8110 15930 8350 16170
rect 8440 15930 8680 16170
rect 8770 15930 9010 16170
rect 9100 15930 9340 16170
rect 9430 15930 9670 16170
rect 9760 15930 10000 16170
rect 10090 15930 10330 16170
rect 10420 15930 10660 16170
rect 10750 15930 10990 16170
rect 11080 15930 11320 16170
rect 11410 15930 11650 16170
rect 11740 15930 11980 16170
rect 12070 15930 12310 16170
rect 12400 15930 12640 16170
rect 12730 15930 12970 16170
rect 13060 15930 13300 16170
rect 13390 15930 13630 16170
rect 13720 15930 13960 16170
rect 14050 15930 14290 16170
rect 14380 15930 14620 16170
rect 14710 15930 14950 16170
rect 15040 15930 15280 16170
rect 15370 15930 15610 16170
rect 15700 15930 15940 16170
rect 16030 15930 16270 16170
rect 16360 15930 16600 16170
rect 16690 15930 16930 16170
rect 17020 15930 17260 16170
rect 17350 15930 17590 16170
rect 17680 15930 17920 16170
rect 18010 15930 18250 16170
rect 18340 15930 18580 16170
rect 18670 15930 18910 16170
rect 19000 15930 19240 16170
rect 19330 15930 19570 16170
rect 7780 15600 8020 15840
rect 8110 15600 8350 15840
rect 8440 15600 8680 15840
rect 8770 15600 9010 15840
rect 9100 15600 9340 15840
rect 9430 15600 9670 15840
rect 9760 15600 10000 15840
rect 10090 15600 10330 15840
rect 10420 15600 10660 15840
rect 10750 15600 10990 15840
rect 11080 15600 11320 15840
rect 11410 15600 11650 15840
rect 11740 15600 11980 15840
rect 12070 15600 12310 15840
rect 12400 15600 12640 15840
rect 12730 15600 12970 15840
rect 13060 15600 13300 15840
rect 13390 15600 13630 15840
rect 13720 15600 13960 15840
rect 14050 15600 14290 15840
rect 14380 15600 14620 15840
rect 14710 15600 14950 15840
rect 15040 15600 15280 15840
rect 15370 15600 15610 15840
rect 15700 15600 15940 15840
rect 16030 15600 16270 15840
rect 16360 15600 16600 15840
rect 16690 15600 16930 15840
rect 17020 15600 17260 15840
rect 17350 15600 17590 15840
rect 17680 15600 17920 15840
rect 18010 15600 18250 15840
rect 18340 15600 18580 15840
rect 18670 15600 18910 15840
rect 19000 15600 19240 15840
rect 19330 15600 19570 15840
rect 7780 15270 8020 15510
rect 8110 15270 8350 15510
rect 8440 15270 8680 15510
rect 8770 15270 9010 15510
rect 9100 15270 9340 15510
rect 9430 15270 9670 15510
rect 9760 15270 10000 15510
rect 10090 15270 10330 15510
rect 10420 15270 10660 15510
rect 10750 15270 10990 15510
rect 11080 15270 11320 15510
rect 11410 15270 11650 15510
rect 11740 15270 11980 15510
rect 12070 15270 12310 15510
rect 12400 15270 12640 15510
rect 12730 15270 12970 15510
rect 13060 15270 13300 15510
rect 13390 15270 13630 15510
rect 13720 15270 13960 15510
rect 14050 15270 14290 15510
rect 14380 15270 14620 15510
rect 14710 15270 14950 15510
rect 15040 15270 15280 15510
rect 15370 15270 15610 15510
rect 15700 15270 15940 15510
rect 16030 15270 16270 15510
rect 16360 15270 16600 15510
rect 16690 15270 16930 15510
rect 17020 15270 17260 15510
rect 17350 15270 17590 15510
rect 17680 15270 17920 15510
rect 18010 15270 18250 15510
rect 18340 15270 18580 15510
rect 18670 15270 18910 15510
rect 19000 15270 19240 15510
rect 19330 15270 19570 15510
rect 7780 14940 8020 15180
rect 8110 14940 8350 15180
rect 8440 14940 8680 15180
rect 8770 14940 9010 15180
rect 9100 14940 9340 15180
rect 9430 14940 9670 15180
rect 9760 14940 10000 15180
rect 10090 14940 10330 15180
rect 10420 14940 10660 15180
rect 10750 14940 10990 15180
rect 11080 14940 11320 15180
rect 11410 14940 11650 15180
rect 11740 14940 11980 15180
rect 12070 14940 12310 15180
rect 12400 14940 12640 15180
rect 12730 14940 12970 15180
rect 13060 14940 13300 15180
rect 13390 14940 13630 15180
rect 13720 14940 13960 15180
rect 14050 14940 14290 15180
rect 14380 14940 14620 15180
rect 14710 14940 14950 15180
rect 15040 14940 15280 15180
rect 15370 14940 15610 15180
rect 15700 14940 15940 15180
rect 16030 14940 16270 15180
rect 16360 14940 16600 15180
rect 16690 14940 16930 15180
rect 17020 14940 17260 15180
rect 17350 14940 17590 15180
rect 17680 14940 17920 15180
rect 18010 14940 18250 15180
rect 18340 14940 18580 15180
rect 18670 14940 18910 15180
rect 19000 14940 19240 15180
rect 19330 14940 19570 15180
rect 7780 14610 8020 14850
rect 8110 14610 8350 14850
rect 8440 14610 8680 14850
rect 8770 14610 9010 14850
rect 9100 14610 9340 14850
rect 9430 14610 9670 14850
rect 9760 14610 10000 14850
rect 10090 14610 10330 14850
rect 10420 14610 10660 14850
rect 10750 14610 10990 14850
rect 11080 14610 11320 14850
rect 11410 14610 11650 14850
rect 11740 14610 11980 14850
rect 12070 14610 12310 14850
rect 12400 14610 12640 14850
rect 12730 14610 12970 14850
rect 13060 14610 13300 14850
rect 13390 14610 13630 14850
rect 13720 14610 13960 14850
rect 14050 14610 14290 14850
rect 14380 14610 14620 14850
rect 14710 14610 14950 14850
rect 15040 14610 15280 14850
rect 15370 14610 15610 14850
rect 15700 14610 15940 14850
rect 16030 14610 16270 14850
rect 16360 14610 16600 14850
rect 16690 14610 16930 14850
rect 17020 14610 17260 14850
rect 17350 14610 17590 14850
rect 17680 14610 17920 14850
rect 18010 14610 18250 14850
rect 18340 14610 18580 14850
rect 18670 14610 18910 14850
rect 19000 14610 19240 14850
rect 19330 14610 19570 14850
rect 7780 14280 8020 14520
rect 8110 14280 8350 14520
rect 8440 14280 8680 14520
rect 8770 14280 9010 14520
rect 9100 14280 9340 14520
rect 9430 14280 9670 14520
rect 9760 14280 10000 14520
rect 10090 14280 10330 14520
rect 10420 14280 10660 14520
rect 10750 14280 10990 14520
rect 11080 14280 11320 14520
rect 11410 14280 11650 14520
rect 11740 14280 11980 14520
rect 12070 14280 12310 14520
rect 12400 14280 12640 14520
rect 12730 14280 12970 14520
rect 13060 14280 13300 14520
rect 13390 14280 13630 14520
rect 13720 14280 13960 14520
rect 14050 14280 14290 14520
rect 14380 14280 14620 14520
rect 14710 14280 14950 14520
rect 15040 14280 15280 14520
rect 15370 14280 15610 14520
rect 15700 14280 15940 14520
rect 16030 14280 16270 14520
rect 16360 14280 16600 14520
rect 16690 14280 16930 14520
rect 17020 14280 17260 14520
rect 17350 14280 17590 14520
rect 17680 14280 17920 14520
rect 18010 14280 18250 14520
rect 18340 14280 18580 14520
rect 18670 14280 18910 14520
rect 19000 14280 19240 14520
rect 19330 14280 19570 14520
rect 7780 13950 8020 14190
rect 8110 13950 8350 14190
rect 8440 13950 8680 14190
rect 8770 13950 9010 14190
rect 9100 13950 9340 14190
rect 9430 13950 9670 14190
rect 9760 13950 10000 14190
rect 10090 13950 10330 14190
rect 10420 13950 10660 14190
rect 10750 13950 10990 14190
rect 11080 13950 11320 14190
rect 11410 13950 11650 14190
rect 11740 13950 11980 14190
rect 12070 13950 12310 14190
rect 12400 13950 12640 14190
rect 12730 13950 12970 14190
rect 13060 13950 13300 14190
rect 13390 13950 13630 14190
rect 13720 13950 13960 14190
rect 14050 13950 14290 14190
rect 14380 13950 14620 14190
rect 14710 13950 14950 14190
rect 15040 13950 15280 14190
rect 15370 13950 15610 14190
rect 15700 13950 15940 14190
rect 16030 13950 16270 14190
rect 16360 13950 16600 14190
rect 16690 13950 16930 14190
rect 17020 13950 17260 14190
rect 17350 13950 17590 14190
rect 17680 13950 17920 14190
rect 18010 13950 18250 14190
rect 18340 13950 18580 14190
rect 18670 13950 18910 14190
rect 19000 13950 19240 14190
rect 19330 13950 19570 14190
rect 7780 13620 8020 13860
rect 8110 13620 8350 13860
rect 8440 13620 8680 13860
rect 8770 13620 9010 13860
rect 9100 13620 9340 13860
rect 9430 13620 9670 13860
rect 9760 13620 10000 13860
rect 10090 13620 10330 13860
rect 10420 13620 10660 13860
rect 10750 13620 10990 13860
rect 11080 13620 11320 13860
rect 11410 13620 11650 13860
rect 11740 13620 11980 13860
rect 12070 13620 12310 13860
rect 12400 13620 12640 13860
rect 12730 13620 12970 13860
rect 13060 13620 13300 13860
rect 13390 13620 13630 13860
rect 13720 13620 13960 13860
rect 14050 13620 14290 13860
rect 14380 13620 14620 13860
rect 14710 13620 14950 13860
rect 15040 13620 15280 13860
rect 15370 13620 15610 13860
rect 15700 13620 15940 13860
rect 16030 13620 16270 13860
rect 16360 13620 16600 13860
rect 16690 13620 16930 13860
rect 17020 13620 17260 13860
rect 17350 13620 17590 13860
rect 17680 13620 17920 13860
rect 18010 13620 18250 13860
rect 18340 13620 18580 13860
rect 18670 13620 18910 13860
rect 19000 13620 19240 13860
rect 19330 13620 19570 13860
rect 7780 13290 8020 13530
rect 8110 13290 8350 13530
rect 8440 13290 8680 13530
rect 8770 13290 9010 13530
rect 9100 13290 9340 13530
rect 9430 13290 9670 13530
rect 9760 13290 10000 13530
rect 10090 13290 10330 13530
rect 10420 13290 10660 13530
rect 10750 13290 10990 13530
rect 11080 13290 11320 13530
rect 11410 13290 11650 13530
rect 11740 13290 11980 13530
rect 12070 13290 12310 13530
rect 12400 13290 12640 13530
rect 12730 13290 12970 13530
rect 13060 13290 13300 13530
rect 13390 13290 13630 13530
rect 13720 13290 13960 13530
rect 14050 13290 14290 13530
rect 14380 13290 14620 13530
rect 14710 13290 14950 13530
rect 15040 13290 15280 13530
rect 15370 13290 15610 13530
rect 15700 13290 15940 13530
rect 16030 13290 16270 13530
rect 16360 13290 16600 13530
rect 16690 13290 16930 13530
rect 17020 13290 17260 13530
rect 17350 13290 17590 13530
rect 17680 13290 17920 13530
rect 18010 13290 18250 13530
rect 18340 13290 18580 13530
rect 18670 13290 18910 13530
rect 19000 13290 19240 13530
rect 19330 13290 19570 13530
rect 7780 12960 8020 13200
rect 8110 12960 8350 13200
rect 8440 12960 8680 13200
rect 8770 12960 9010 13200
rect 9100 12960 9340 13200
rect 9430 12960 9670 13200
rect 9760 12960 10000 13200
rect 10090 12960 10330 13200
rect 10420 12960 10660 13200
rect 10750 12960 10990 13200
rect 11080 12960 11320 13200
rect 11410 12960 11650 13200
rect 11740 12960 11980 13200
rect 12070 12960 12310 13200
rect 12400 12960 12640 13200
rect 12730 12960 12970 13200
rect 13060 12960 13300 13200
rect 13390 12960 13630 13200
rect 13720 12960 13960 13200
rect 14050 12960 14290 13200
rect 14380 12960 14620 13200
rect 14710 12960 14950 13200
rect 15040 12960 15280 13200
rect 15370 12960 15610 13200
rect 15700 12960 15940 13200
rect 16030 12960 16270 13200
rect 16360 12960 16600 13200
rect 16690 12960 16930 13200
rect 17020 12960 17260 13200
rect 17350 12960 17590 13200
rect 17680 12960 17920 13200
rect 18010 12960 18250 13200
rect 18340 12960 18580 13200
rect 18670 12960 18910 13200
rect 19000 12960 19240 13200
rect 19330 12960 19570 13200
rect 7780 12630 8020 12870
rect 8110 12630 8350 12870
rect 8440 12630 8680 12870
rect 8770 12630 9010 12870
rect 9100 12630 9340 12870
rect 9430 12630 9670 12870
rect 9760 12630 10000 12870
rect 10090 12630 10330 12870
rect 10420 12630 10660 12870
rect 10750 12630 10990 12870
rect 11080 12630 11320 12870
rect 11410 12630 11650 12870
rect 11740 12630 11980 12870
rect 12070 12630 12310 12870
rect 12400 12630 12640 12870
rect 12730 12630 12970 12870
rect 13060 12630 13300 12870
rect 13390 12630 13630 12870
rect 13720 12630 13960 12870
rect 14050 12630 14290 12870
rect 14380 12630 14620 12870
rect 14710 12630 14950 12870
rect 15040 12630 15280 12870
rect 15370 12630 15610 12870
rect 15700 12630 15940 12870
rect 16030 12630 16270 12870
rect 16360 12630 16600 12870
rect 16690 12630 16930 12870
rect 17020 12630 17260 12870
rect 17350 12630 17590 12870
rect 17680 12630 17920 12870
rect 18010 12630 18250 12870
rect 18340 12630 18580 12870
rect 18670 12630 18910 12870
rect 19000 12630 19240 12870
rect 19330 12630 19570 12870
rect 7780 12300 8020 12540
rect 8110 12300 8350 12540
rect 8440 12300 8680 12540
rect 8770 12300 9010 12540
rect 9100 12300 9340 12540
rect 9430 12300 9670 12540
rect 9760 12300 10000 12540
rect 10090 12300 10330 12540
rect 10420 12300 10660 12540
rect 10750 12300 10990 12540
rect 11080 12300 11320 12540
rect 11410 12300 11650 12540
rect 11740 12300 11980 12540
rect 12070 12300 12310 12540
rect 12400 12300 12640 12540
rect 12730 12300 12970 12540
rect 13060 12300 13300 12540
rect 13390 12300 13630 12540
rect 13720 12300 13960 12540
rect 14050 12300 14290 12540
rect 14380 12300 14620 12540
rect 14710 12300 14950 12540
rect 15040 12300 15280 12540
rect 15370 12300 15610 12540
rect 15700 12300 15940 12540
rect 16030 12300 16270 12540
rect 16360 12300 16600 12540
rect 16690 12300 16930 12540
rect 17020 12300 17260 12540
rect 17350 12300 17590 12540
rect 17680 12300 17920 12540
rect 18010 12300 18250 12540
rect 18340 12300 18580 12540
rect 18670 12300 18910 12540
rect 19000 12300 19240 12540
rect 19330 12300 19570 12540
rect 7780 11970 8020 12210
rect 8110 11970 8350 12210
rect 8440 11970 8680 12210
rect 8770 11970 9010 12210
rect 9100 11970 9340 12210
rect 9430 11970 9670 12210
rect 9760 11970 10000 12210
rect 10090 11970 10330 12210
rect 10420 11970 10660 12210
rect 10750 11970 10990 12210
rect 11080 11970 11320 12210
rect 11410 11970 11650 12210
rect 11740 11970 11980 12210
rect 12070 11970 12310 12210
rect 12400 11970 12640 12210
rect 12730 11970 12970 12210
rect 13060 11970 13300 12210
rect 13390 11970 13630 12210
rect 13720 11970 13960 12210
rect 14050 11970 14290 12210
rect 14380 11970 14620 12210
rect 14710 11970 14950 12210
rect 15040 11970 15280 12210
rect 15370 11970 15610 12210
rect 15700 11970 15940 12210
rect 16030 11970 16270 12210
rect 16360 11970 16600 12210
rect 16690 11970 16930 12210
rect 17020 11970 17260 12210
rect 17350 11970 17590 12210
rect 17680 11970 17920 12210
rect 18010 11970 18250 12210
rect 18340 11970 18580 12210
rect 18670 11970 18910 12210
rect 19000 11970 19240 12210
rect 19330 11970 19570 12210
rect 7780 11640 8020 11880
rect 8110 11640 8350 11880
rect 8440 11640 8680 11880
rect 8770 11640 9010 11880
rect 9100 11640 9340 11880
rect 9430 11640 9670 11880
rect 9760 11640 10000 11880
rect 10090 11640 10330 11880
rect 10420 11640 10660 11880
rect 10750 11640 10990 11880
rect 11080 11640 11320 11880
rect 11410 11640 11650 11880
rect 11740 11640 11980 11880
rect 12070 11640 12310 11880
rect 12400 11640 12640 11880
rect 12730 11640 12970 11880
rect 13060 11640 13300 11880
rect 13390 11640 13630 11880
rect 13720 11640 13960 11880
rect 14050 11640 14290 11880
rect 14380 11640 14620 11880
rect 14710 11640 14950 11880
rect 15040 11640 15280 11880
rect 15370 11640 15610 11880
rect 15700 11640 15940 11880
rect 16030 11640 16270 11880
rect 16360 11640 16600 11880
rect 16690 11640 16930 11880
rect 17020 11640 17260 11880
rect 17350 11640 17590 11880
rect 17680 11640 17920 11880
rect 18010 11640 18250 11880
rect 18340 11640 18580 11880
rect 18670 11640 18910 11880
rect 19000 11640 19240 11880
rect 19330 11640 19570 11880
rect 7780 11310 8020 11550
rect 8110 11310 8350 11550
rect 8440 11310 8680 11550
rect 8770 11310 9010 11550
rect 9100 11310 9340 11550
rect 9430 11310 9670 11550
rect 9760 11310 10000 11550
rect 10090 11310 10330 11550
rect 10420 11310 10660 11550
rect 10750 11310 10990 11550
rect 11080 11310 11320 11550
rect 11410 11310 11650 11550
rect 11740 11310 11980 11550
rect 12070 11310 12310 11550
rect 12400 11310 12640 11550
rect 12730 11310 12970 11550
rect 13060 11310 13300 11550
rect 13390 11310 13630 11550
rect 13720 11310 13960 11550
rect 14050 11310 14290 11550
rect 14380 11310 14620 11550
rect 14710 11310 14950 11550
rect 15040 11310 15280 11550
rect 15370 11310 15610 11550
rect 15700 11310 15940 11550
rect 16030 11310 16270 11550
rect 16360 11310 16600 11550
rect 16690 11310 16930 11550
rect 17020 11310 17260 11550
rect 17350 11310 17590 11550
rect 17680 11310 17920 11550
rect 18010 11310 18250 11550
rect 18340 11310 18580 11550
rect 18670 11310 18910 11550
rect 19000 11310 19240 11550
rect 19330 11310 19570 11550
rect 7780 10980 8020 11220
rect 8110 10980 8350 11220
rect 8440 10980 8680 11220
rect 8770 10980 9010 11220
rect 9100 10980 9340 11220
rect 9430 10980 9670 11220
rect 9760 10980 10000 11220
rect 10090 10980 10330 11220
rect 10420 10980 10660 11220
rect 10750 10980 10990 11220
rect 11080 10980 11320 11220
rect 11410 10980 11650 11220
rect 11740 10980 11980 11220
rect 12070 10980 12310 11220
rect 12400 10980 12640 11220
rect 12730 10980 12970 11220
rect 13060 10980 13300 11220
rect 13390 10980 13630 11220
rect 13720 10980 13960 11220
rect 14050 10980 14290 11220
rect 14380 10980 14620 11220
rect 14710 10980 14950 11220
rect 15040 10980 15280 11220
rect 15370 10980 15610 11220
rect 15700 10980 15940 11220
rect 16030 10980 16270 11220
rect 16360 10980 16600 11220
rect 16690 10980 16930 11220
rect 17020 10980 17260 11220
rect 17350 10980 17590 11220
rect 17680 10980 17920 11220
rect 18010 10980 18250 11220
rect 18340 10980 18580 11220
rect 18670 10980 18910 11220
rect 19000 10980 19240 11220
rect 19330 10980 19570 11220
rect 7780 10650 8020 10890
rect 8110 10650 8350 10890
rect 8440 10650 8680 10890
rect 8770 10650 9010 10890
rect 9100 10650 9340 10890
rect 9430 10650 9670 10890
rect 9760 10650 10000 10890
rect 10090 10650 10330 10890
rect 10420 10650 10660 10890
rect 10750 10650 10990 10890
rect 11080 10650 11320 10890
rect 11410 10650 11650 10890
rect 11740 10650 11980 10890
rect 12070 10650 12310 10890
rect 12400 10650 12640 10890
rect 12730 10650 12970 10890
rect 13060 10650 13300 10890
rect 13390 10650 13630 10890
rect 13720 10650 13960 10890
rect 14050 10650 14290 10890
rect 14380 10650 14620 10890
rect 14710 10650 14950 10890
rect 15040 10650 15280 10890
rect 15370 10650 15610 10890
rect 15700 10650 15940 10890
rect 16030 10650 16270 10890
rect 16360 10650 16600 10890
rect 16690 10650 16930 10890
rect 17020 10650 17260 10890
rect 17350 10650 17590 10890
rect 17680 10650 17920 10890
rect 18010 10650 18250 10890
rect 18340 10650 18580 10890
rect 18670 10650 18910 10890
rect 19000 10650 19240 10890
rect 19330 10650 19570 10890
rect 7780 10320 8020 10560
rect 8110 10320 8350 10560
rect 8440 10320 8680 10560
rect 8770 10320 9010 10560
rect 9100 10320 9340 10560
rect 9430 10320 9670 10560
rect 9760 10320 10000 10560
rect 10090 10320 10330 10560
rect 10420 10320 10660 10560
rect 10750 10320 10990 10560
rect 11080 10320 11320 10560
rect 11410 10320 11650 10560
rect 11740 10320 11980 10560
rect 12070 10320 12310 10560
rect 12400 10320 12640 10560
rect 12730 10320 12970 10560
rect 13060 10320 13300 10560
rect 13390 10320 13630 10560
rect 13720 10320 13960 10560
rect 14050 10320 14290 10560
rect 14380 10320 14620 10560
rect 14710 10320 14950 10560
rect 15040 10320 15280 10560
rect 15370 10320 15610 10560
rect 15700 10320 15940 10560
rect 16030 10320 16270 10560
rect 16360 10320 16600 10560
rect 16690 10320 16930 10560
rect 17020 10320 17260 10560
rect 17350 10320 17590 10560
rect 17680 10320 17920 10560
rect 18010 10320 18250 10560
rect 18340 10320 18580 10560
rect 18670 10320 18910 10560
rect 19000 10320 19240 10560
rect 19330 10320 19570 10560
rect 7780 9990 8020 10230
rect 8110 9990 8350 10230
rect 8440 9990 8680 10230
rect 8770 9990 9010 10230
rect 9100 9990 9340 10230
rect 9430 9990 9670 10230
rect 9760 9990 10000 10230
rect 10090 9990 10330 10230
rect 10420 9990 10660 10230
rect 10750 9990 10990 10230
rect 11080 9990 11320 10230
rect 11410 9990 11650 10230
rect 11740 9990 11980 10230
rect 12070 9990 12310 10230
rect 12400 9990 12640 10230
rect 12730 9990 12970 10230
rect 13060 9990 13300 10230
rect 13390 9990 13630 10230
rect 13720 9990 13960 10230
rect 14050 9990 14290 10230
rect 14380 9990 14620 10230
rect 14710 9990 14950 10230
rect 15040 9990 15280 10230
rect 15370 9990 15610 10230
rect 15700 9990 15940 10230
rect 16030 9990 16270 10230
rect 16360 9990 16600 10230
rect 16690 9990 16930 10230
rect 17020 9990 17260 10230
rect 17350 9990 17590 10230
rect 17680 9990 17920 10230
rect 18010 9990 18250 10230
rect 18340 9990 18580 10230
rect 18670 9990 18910 10230
rect 19000 9990 19240 10230
rect 19330 9990 19570 10230
rect 7780 9660 8020 9900
rect 8110 9660 8350 9900
rect 8440 9660 8680 9900
rect 8770 9660 9010 9900
rect 9100 9660 9340 9900
rect 9430 9660 9670 9900
rect 9760 9660 10000 9900
rect 10090 9660 10330 9900
rect 10420 9660 10660 9900
rect 10750 9660 10990 9900
rect 11080 9660 11320 9900
rect 11410 9660 11650 9900
rect 11740 9660 11980 9900
rect 12070 9660 12310 9900
rect 12400 9660 12640 9900
rect 12730 9660 12970 9900
rect 13060 9660 13300 9900
rect 13390 9660 13630 9900
rect 13720 9660 13960 9900
rect 14050 9660 14290 9900
rect 14380 9660 14620 9900
rect 14710 9660 14950 9900
rect 15040 9660 15280 9900
rect 15370 9660 15610 9900
rect 15700 9660 15940 9900
rect 16030 9660 16270 9900
rect 16360 9660 16600 9900
rect 16690 9660 16930 9900
rect 17020 9660 17260 9900
rect 17350 9660 17590 9900
rect 17680 9660 17920 9900
rect 18010 9660 18250 9900
rect 18340 9660 18580 9900
rect 18670 9660 18910 9900
rect 19000 9660 19240 9900
rect 19330 9660 19570 9900
rect 7780 9330 8020 9570
rect 8110 9330 8350 9570
rect 8440 9330 8680 9570
rect 8770 9330 9010 9570
rect 9100 9330 9340 9570
rect 9430 9330 9670 9570
rect 9760 9330 10000 9570
rect 10090 9330 10330 9570
rect 10420 9330 10660 9570
rect 10750 9330 10990 9570
rect 11080 9330 11320 9570
rect 11410 9330 11650 9570
rect 11740 9330 11980 9570
rect 12070 9330 12310 9570
rect 12400 9330 12640 9570
rect 12730 9330 12970 9570
rect 13060 9330 13300 9570
rect 13390 9330 13630 9570
rect 13720 9330 13960 9570
rect 14050 9330 14290 9570
rect 14380 9330 14620 9570
rect 14710 9330 14950 9570
rect 15040 9330 15280 9570
rect 15370 9330 15610 9570
rect 15700 9330 15940 9570
rect 16030 9330 16270 9570
rect 16360 9330 16600 9570
rect 16690 9330 16930 9570
rect 17020 9330 17260 9570
rect 17350 9330 17590 9570
rect 17680 9330 17920 9570
rect 18010 9330 18250 9570
rect 18340 9330 18580 9570
rect 18670 9330 18910 9570
rect 19000 9330 19240 9570
rect 19330 9330 19570 9570
rect 7780 9000 8020 9240
rect 8110 9000 8350 9240
rect 8440 9000 8680 9240
rect 8770 9000 9010 9240
rect 9100 9000 9340 9240
rect 9430 9000 9670 9240
rect 9760 9000 10000 9240
rect 10090 9000 10330 9240
rect 10420 9000 10660 9240
rect 10750 9000 10990 9240
rect 11080 9000 11320 9240
rect 11410 9000 11650 9240
rect 11740 9000 11980 9240
rect 12070 9000 12310 9240
rect 12400 9000 12640 9240
rect 12730 9000 12970 9240
rect 13060 9000 13300 9240
rect 13390 9000 13630 9240
rect 13720 9000 13960 9240
rect 14050 9000 14290 9240
rect 14380 9000 14620 9240
rect 14710 9000 14950 9240
rect 15040 9000 15280 9240
rect 15370 9000 15610 9240
rect 15700 9000 15940 9240
rect 16030 9000 16270 9240
rect 16360 9000 16600 9240
rect 16690 9000 16930 9240
rect 17020 9000 17260 9240
rect 17350 9000 17590 9240
rect 17680 9000 17920 9240
rect 18010 9000 18250 9240
rect 18340 9000 18580 9240
rect 18670 9000 18910 9240
rect 19000 9000 19240 9240
rect 19330 9000 19570 9240
rect 28780 7590 29020 7830
rect 29110 7590 29350 7830
rect 29440 7590 29680 7830
rect 29770 7590 30010 7830
rect 30100 7590 30340 7830
rect 30430 7590 30670 7830
rect 30760 7590 31000 7830
rect 31090 7590 31330 7830
rect 31420 7590 31660 7830
rect 31750 7590 31990 7830
rect 32080 7590 32320 7830
rect 32410 7590 32650 7830
rect 32740 7590 32980 7830
rect 33070 7590 33310 7830
rect 33400 7590 33640 7830
rect 33730 7590 33970 7830
rect 34060 7590 34300 7830
rect 34390 7590 34630 7830
rect 34720 7590 34960 7830
rect 35050 7590 35290 7830
rect 28780 7260 29020 7500
rect 29110 7260 29350 7500
rect 29440 7260 29680 7500
rect 29770 7260 30010 7500
rect 30100 7260 30340 7500
rect 30430 7260 30670 7500
rect 30760 7260 31000 7500
rect 31090 7260 31330 7500
rect 31420 7260 31660 7500
rect 31750 7260 31990 7500
rect 32080 7260 32320 7500
rect 32410 7260 32650 7500
rect 32740 7260 32980 7500
rect 33070 7260 33310 7500
rect 33400 7260 33640 7500
rect 33730 7260 33970 7500
rect 34060 7260 34300 7500
rect 34390 7260 34630 7500
rect 34720 7260 34960 7500
rect 35050 7260 35290 7500
rect 28780 6930 29020 7170
rect 29110 6930 29350 7170
rect 29440 6930 29680 7170
rect 29770 6930 30010 7170
rect 30100 6930 30340 7170
rect 30430 6930 30670 7170
rect 30760 6930 31000 7170
rect 31090 6930 31330 7170
rect 31420 6930 31660 7170
rect 31750 6930 31990 7170
rect 32080 6930 32320 7170
rect 32410 6930 32650 7170
rect 32740 6930 32980 7170
rect 33070 6930 33310 7170
rect 33400 6930 33640 7170
rect 33730 6930 33970 7170
rect 34060 6930 34300 7170
rect 34390 6930 34630 7170
rect 34720 6930 34960 7170
rect 35050 6930 35290 7170
rect 28780 6600 29020 6840
rect 29110 6600 29350 6840
rect 29440 6600 29680 6840
rect 29770 6600 30010 6840
rect 30100 6600 30340 6840
rect 30430 6600 30670 6840
rect 30760 6600 31000 6840
rect 31090 6600 31330 6840
rect 31420 6600 31660 6840
rect 31750 6600 31990 6840
rect 32080 6600 32320 6840
rect 32410 6600 32650 6840
rect 32740 6600 32980 6840
rect 33070 6600 33310 6840
rect 33400 6600 33640 6840
rect 33730 6600 33970 6840
rect 34060 6600 34300 6840
rect 34390 6600 34630 6840
rect 34720 6600 34960 6840
rect 35050 6600 35290 6840
rect 28780 6270 29020 6510
rect 29110 6270 29350 6510
rect 29440 6270 29680 6510
rect 29770 6270 30010 6510
rect 30100 6270 30340 6510
rect 30430 6270 30670 6510
rect 30760 6270 31000 6510
rect 31090 6270 31330 6510
rect 31420 6270 31660 6510
rect 31750 6270 31990 6510
rect 32080 6270 32320 6510
rect 32410 6270 32650 6510
rect 32740 6270 32980 6510
rect 33070 6270 33310 6510
rect 33400 6270 33640 6510
rect 33730 6270 33970 6510
rect 34060 6270 34300 6510
rect 34390 6270 34630 6510
rect 34720 6270 34960 6510
rect 35050 6270 35290 6510
rect 28780 5940 29020 6180
rect 29110 5940 29350 6180
rect 29440 5940 29680 6180
rect 29770 5940 30010 6180
rect 30100 5940 30340 6180
rect 30430 5940 30670 6180
rect 30760 5940 31000 6180
rect 31090 5940 31330 6180
rect 31420 5940 31660 6180
rect 31750 5940 31990 6180
rect 32080 5940 32320 6180
rect 32410 5940 32650 6180
rect 32740 5940 32980 6180
rect 33070 5940 33310 6180
rect 33400 5940 33640 6180
rect 33730 5940 33970 6180
rect 34060 5940 34300 6180
rect 34390 5940 34630 6180
rect 34720 5940 34960 6180
rect 35050 5940 35290 6180
rect 28780 5610 29020 5850
rect 29110 5610 29350 5850
rect 29440 5610 29680 5850
rect 29770 5610 30010 5850
rect 30100 5610 30340 5850
rect 30430 5610 30670 5850
rect 30760 5610 31000 5850
rect 31090 5610 31330 5850
rect 31420 5610 31660 5850
rect 31750 5610 31990 5850
rect 32080 5610 32320 5850
rect 32410 5610 32650 5850
rect 32740 5610 32980 5850
rect 33070 5610 33310 5850
rect 33400 5610 33640 5850
rect 33730 5610 33970 5850
rect 34060 5610 34300 5850
rect 34390 5610 34630 5850
rect 34720 5610 34960 5850
rect 35050 5610 35290 5850
rect 28780 5280 29020 5520
rect 29110 5280 29350 5520
rect 29440 5280 29680 5520
rect 29770 5280 30010 5520
rect 30100 5280 30340 5520
rect 30430 5280 30670 5520
rect 30760 5280 31000 5520
rect 31090 5280 31330 5520
rect 31420 5280 31660 5520
rect 31750 5280 31990 5520
rect 32080 5280 32320 5520
rect 32410 5280 32650 5520
rect 32740 5280 32980 5520
rect 33070 5280 33310 5520
rect 33400 5280 33640 5520
rect 33730 5280 33970 5520
rect 34060 5280 34300 5520
rect 34390 5280 34630 5520
rect 34720 5280 34960 5520
rect 35050 5280 35290 5520
rect 28780 4950 29020 5190
rect 29110 4950 29350 5190
rect 29440 4950 29680 5190
rect 29770 4950 30010 5190
rect 30100 4950 30340 5190
rect 30430 4950 30670 5190
rect 30760 4950 31000 5190
rect 31090 4950 31330 5190
rect 31420 4950 31660 5190
rect 31750 4950 31990 5190
rect 32080 4950 32320 5190
rect 32410 4950 32650 5190
rect 32740 4950 32980 5190
rect 33070 4950 33310 5190
rect 33400 4950 33640 5190
rect 33730 4950 33970 5190
rect 34060 4950 34300 5190
rect 34390 4950 34630 5190
rect 34720 4950 34960 5190
rect 35050 4950 35290 5190
rect 28780 4620 29020 4860
rect 29110 4620 29350 4860
rect 29440 4620 29680 4860
rect 29770 4620 30010 4860
rect 30100 4620 30340 4860
rect 30430 4620 30670 4860
rect 30760 4620 31000 4860
rect 31090 4620 31330 4860
rect 31420 4620 31660 4860
rect 31750 4620 31990 4860
rect 32080 4620 32320 4860
rect 32410 4620 32650 4860
rect 32740 4620 32980 4860
rect 33070 4620 33310 4860
rect 33400 4620 33640 4860
rect 33730 4620 33970 4860
rect 34060 4620 34300 4860
rect 34390 4620 34630 4860
rect 34720 4620 34960 4860
rect 35050 4620 35290 4860
rect 28780 4290 29020 4530
rect 29110 4290 29350 4530
rect 29440 4290 29680 4530
rect 29770 4290 30010 4530
rect 30100 4290 30340 4530
rect 30430 4290 30670 4530
rect 30760 4290 31000 4530
rect 31090 4290 31330 4530
rect 31420 4290 31660 4530
rect 31750 4290 31990 4530
rect 32080 4290 32320 4530
rect 32410 4290 32650 4530
rect 32740 4290 32980 4530
rect 33070 4290 33310 4530
rect 33400 4290 33640 4530
rect 33730 4290 33970 4530
rect 34060 4290 34300 4530
rect 34390 4290 34630 4530
rect 34720 4290 34960 4530
rect 35050 4290 35290 4530
rect 28780 3960 29020 4200
rect 29110 3960 29350 4200
rect 29440 3960 29680 4200
rect 29770 3960 30010 4200
rect 30100 3960 30340 4200
rect 30430 3960 30670 4200
rect 30760 3960 31000 4200
rect 31090 3960 31330 4200
rect 31420 3960 31660 4200
rect 31750 3960 31990 4200
rect 32080 3960 32320 4200
rect 32410 3960 32650 4200
rect 32740 3960 32980 4200
rect 33070 3960 33310 4200
rect 33400 3960 33640 4200
rect 33730 3960 33970 4200
rect 34060 3960 34300 4200
rect 34390 3960 34630 4200
rect 34720 3960 34960 4200
rect 35050 3960 35290 4200
rect 28780 3630 29020 3870
rect 29110 3630 29350 3870
rect 29440 3630 29680 3870
rect 29770 3630 30010 3870
rect 30100 3630 30340 3870
rect 30430 3630 30670 3870
rect 30760 3630 31000 3870
rect 31090 3630 31330 3870
rect 31420 3630 31660 3870
rect 31750 3630 31990 3870
rect 32080 3630 32320 3870
rect 32410 3630 32650 3870
rect 32740 3630 32980 3870
rect 33070 3630 33310 3870
rect 33400 3630 33640 3870
rect 33730 3630 33970 3870
rect 34060 3630 34300 3870
rect 34390 3630 34630 3870
rect 34720 3630 34960 3870
rect 35050 3630 35290 3870
rect 28780 3300 29020 3540
rect 29110 3300 29350 3540
rect 29440 3300 29680 3540
rect 29770 3300 30010 3540
rect 30100 3300 30340 3540
rect 30430 3300 30670 3540
rect 30760 3300 31000 3540
rect 31090 3300 31330 3540
rect 31420 3300 31660 3540
rect 31750 3300 31990 3540
rect 32080 3300 32320 3540
rect 32410 3300 32650 3540
rect 32740 3300 32980 3540
rect 33070 3300 33310 3540
rect 33400 3300 33640 3540
rect 33730 3300 33970 3540
rect 34060 3300 34300 3540
rect 34390 3300 34630 3540
rect 34720 3300 34960 3540
rect 35050 3300 35290 3540
rect 28780 2970 29020 3210
rect 29110 2970 29350 3210
rect 29440 2970 29680 3210
rect 29770 2970 30010 3210
rect 30100 2970 30340 3210
rect 30430 2970 30670 3210
rect 30760 2970 31000 3210
rect 31090 2970 31330 3210
rect 31420 2970 31660 3210
rect 31750 2970 31990 3210
rect 32080 2970 32320 3210
rect 32410 2970 32650 3210
rect 32740 2970 32980 3210
rect 33070 2970 33310 3210
rect 33400 2970 33640 3210
rect 33730 2970 33970 3210
rect 34060 2970 34300 3210
rect 34390 2970 34630 3210
rect 34720 2970 34960 3210
rect 35050 2970 35290 3210
rect 28780 2640 29020 2880
rect 29110 2640 29350 2880
rect 29440 2640 29680 2880
rect 29770 2640 30010 2880
rect 30100 2640 30340 2880
rect 30430 2640 30670 2880
rect 30760 2640 31000 2880
rect 31090 2640 31330 2880
rect 31420 2640 31660 2880
rect 31750 2640 31990 2880
rect 32080 2640 32320 2880
rect 32410 2640 32650 2880
rect 32740 2640 32980 2880
rect 33070 2640 33310 2880
rect 33400 2640 33640 2880
rect 33730 2640 33970 2880
rect 34060 2640 34300 2880
rect 34390 2640 34630 2880
rect 34720 2640 34960 2880
rect 35050 2640 35290 2880
rect 28780 2310 29020 2550
rect 29110 2310 29350 2550
rect 29440 2310 29680 2550
rect 29770 2310 30010 2550
rect 30100 2310 30340 2550
rect 30430 2310 30670 2550
rect 30760 2310 31000 2550
rect 31090 2310 31330 2550
rect 31420 2310 31660 2550
rect 31750 2310 31990 2550
rect 32080 2310 32320 2550
rect 32410 2310 32650 2550
rect 32740 2310 32980 2550
rect 33070 2310 33310 2550
rect 33400 2310 33640 2550
rect 33730 2310 33970 2550
rect 34060 2310 34300 2550
rect 34390 2310 34630 2550
rect 34720 2310 34960 2550
rect 35050 2310 35290 2550
rect 28780 1980 29020 2220
rect 29110 1980 29350 2220
rect 29440 1980 29680 2220
rect 29770 1980 30010 2220
rect 30100 1980 30340 2220
rect 30430 1980 30670 2220
rect 30760 1980 31000 2220
rect 31090 1980 31330 2220
rect 31420 1980 31660 2220
rect 31750 1980 31990 2220
rect 32080 1980 32320 2220
rect 32410 1980 32650 2220
rect 32740 1980 32980 2220
rect 33070 1980 33310 2220
rect 33400 1980 33640 2220
rect 33730 1980 33970 2220
rect 34060 1980 34300 2220
rect 34390 1980 34630 2220
rect 34720 1980 34960 2220
rect 35050 1980 35290 2220
rect 28780 1650 29020 1890
rect 29110 1650 29350 1890
rect 29440 1650 29680 1890
rect 29770 1650 30010 1890
rect 30100 1650 30340 1890
rect 30430 1650 30670 1890
rect 30760 1650 31000 1890
rect 31090 1650 31330 1890
rect 31420 1650 31660 1890
rect 31750 1650 31990 1890
rect 32080 1650 32320 1890
rect 32410 1650 32650 1890
rect 32740 1650 32980 1890
rect 33070 1650 33310 1890
rect 33400 1650 33640 1890
rect 33730 1650 33970 1890
rect 34060 1650 34300 1890
rect 34390 1650 34630 1890
rect 34720 1650 34960 1890
rect 35050 1650 35290 1890
rect 28780 1320 29020 1560
rect 29110 1320 29350 1560
rect 29440 1320 29680 1560
rect 29770 1320 30010 1560
rect 30100 1320 30340 1560
rect 30430 1320 30670 1560
rect 30760 1320 31000 1560
rect 31090 1320 31330 1560
rect 31420 1320 31660 1560
rect 31750 1320 31990 1560
rect 32080 1320 32320 1560
rect 32410 1320 32650 1560
rect 32740 1320 32980 1560
rect 33070 1320 33310 1560
rect 33400 1320 33640 1560
rect 33730 1320 33970 1560
rect 34060 1320 34300 1560
rect 34390 1320 34630 1560
rect 34720 1320 34960 1560
rect 35050 1320 35290 1560
rect 28780 -10 29020 230
rect 29110 -10 29350 230
rect 29440 -10 29680 230
rect 29770 -10 30010 230
rect 30100 -10 30340 230
rect 30430 -10 30670 230
rect 30760 -10 31000 230
rect 31090 -10 31330 230
rect 31420 -10 31660 230
rect 31750 -10 31990 230
rect 32080 -10 32320 230
rect 32410 -10 32650 230
rect 32740 -10 32980 230
rect 33070 -10 33310 230
rect 33400 -10 33640 230
rect 33730 -10 33970 230
rect 34060 -10 34300 230
rect 34390 -10 34630 230
rect 34720 -10 34960 230
rect 35050 -10 35290 230
rect 28780 -340 29020 -100
rect 29110 -340 29350 -100
rect 29440 -340 29680 -100
rect 29770 -340 30010 -100
rect 30100 -340 30340 -100
rect 30430 -340 30670 -100
rect 30760 -340 31000 -100
rect 31090 -340 31330 -100
rect 31420 -340 31660 -100
rect 31750 -340 31990 -100
rect 32080 -340 32320 -100
rect 32410 -340 32650 -100
rect 32740 -340 32980 -100
rect 33070 -340 33310 -100
rect 33400 -340 33640 -100
rect 33730 -340 33970 -100
rect 34060 -340 34300 -100
rect 34390 -340 34630 -100
rect 34720 -340 34960 -100
rect 35050 -340 35290 -100
rect 28780 -670 29020 -430
rect 29110 -670 29350 -430
rect 29440 -670 29680 -430
rect 29770 -670 30010 -430
rect 30100 -670 30340 -430
rect 30430 -670 30670 -430
rect 30760 -670 31000 -430
rect 31090 -670 31330 -430
rect 31420 -670 31660 -430
rect 31750 -670 31990 -430
rect 32080 -670 32320 -430
rect 32410 -670 32650 -430
rect 32740 -670 32980 -430
rect 33070 -670 33310 -430
rect 33400 -670 33640 -430
rect 33730 -670 33970 -430
rect 34060 -670 34300 -430
rect 34390 -670 34630 -430
rect 34720 -670 34960 -430
rect 35050 -670 35290 -430
rect 28780 -1000 29020 -760
rect 29110 -1000 29350 -760
rect 29440 -1000 29680 -760
rect 29770 -1000 30010 -760
rect 30100 -1000 30340 -760
rect 30430 -1000 30670 -760
rect 30760 -1000 31000 -760
rect 31090 -1000 31330 -760
rect 31420 -1000 31660 -760
rect 31750 -1000 31990 -760
rect 32080 -1000 32320 -760
rect 32410 -1000 32650 -760
rect 32740 -1000 32980 -760
rect 33070 -1000 33310 -760
rect 33400 -1000 33640 -760
rect 33730 -1000 33970 -760
rect 34060 -1000 34300 -760
rect 34390 -1000 34630 -760
rect 34720 -1000 34960 -760
rect 35050 -1000 35290 -760
rect 28780 -1330 29020 -1090
rect 29110 -1330 29350 -1090
rect 29440 -1330 29680 -1090
rect 29770 -1330 30010 -1090
rect 30100 -1330 30340 -1090
rect 30430 -1330 30670 -1090
rect 30760 -1330 31000 -1090
rect 31090 -1330 31330 -1090
rect 31420 -1330 31660 -1090
rect 31750 -1330 31990 -1090
rect 32080 -1330 32320 -1090
rect 32410 -1330 32650 -1090
rect 32740 -1330 32980 -1090
rect 33070 -1330 33310 -1090
rect 33400 -1330 33640 -1090
rect 33730 -1330 33970 -1090
rect 34060 -1330 34300 -1090
rect 34390 -1330 34630 -1090
rect 34720 -1330 34960 -1090
rect 35050 -1330 35290 -1090
rect 28780 -1660 29020 -1420
rect 29110 -1660 29350 -1420
rect 29440 -1660 29680 -1420
rect 29770 -1660 30010 -1420
rect 30100 -1660 30340 -1420
rect 30430 -1660 30670 -1420
rect 30760 -1660 31000 -1420
rect 31090 -1660 31330 -1420
rect 31420 -1660 31660 -1420
rect 31750 -1660 31990 -1420
rect 32080 -1660 32320 -1420
rect 32410 -1660 32650 -1420
rect 32740 -1660 32980 -1420
rect 33070 -1660 33310 -1420
rect 33400 -1660 33640 -1420
rect 33730 -1660 33970 -1420
rect 34060 -1660 34300 -1420
rect 34390 -1660 34630 -1420
rect 34720 -1660 34960 -1420
rect 35050 -1660 35290 -1420
rect 28780 -1990 29020 -1750
rect 29110 -1990 29350 -1750
rect 29440 -1990 29680 -1750
rect 29770 -1990 30010 -1750
rect 30100 -1990 30340 -1750
rect 30430 -1990 30670 -1750
rect 30760 -1990 31000 -1750
rect 31090 -1990 31330 -1750
rect 31420 -1990 31660 -1750
rect 31750 -1990 31990 -1750
rect 32080 -1990 32320 -1750
rect 32410 -1990 32650 -1750
rect 32740 -1990 32980 -1750
rect 33070 -1990 33310 -1750
rect 33400 -1990 33640 -1750
rect 33730 -1990 33970 -1750
rect 34060 -1990 34300 -1750
rect 34390 -1990 34630 -1750
rect 34720 -1990 34960 -1750
rect 35050 -1990 35290 -1750
rect 28780 -2320 29020 -2080
rect 29110 -2320 29350 -2080
rect 29440 -2320 29680 -2080
rect 29770 -2320 30010 -2080
rect 30100 -2320 30340 -2080
rect 30430 -2320 30670 -2080
rect 30760 -2320 31000 -2080
rect 31090 -2320 31330 -2080
rect 31420 -2320 31660 -2080
rect 31750 -2320 31990 -2080
rect 32080 -2320 32320 -2080
rect 32410 -2320 32650 -2080
rect 32740 -2320 32980 -2080
rect 33070 -2320 33310 -2080
rect 33400 -2320 33640 -2080
rect 33730 -2320 33970 -2080
rect 34060 -2320 34300 -2080
rect 34390 -2320 34630 -2080
rect 34720 -2320 34960 -2080
rect 35050 -2320 35290 -2080
rect 28780 -2650 29020 -2410
rect 29110 -2650 29350 -2410
rect 29440 -2650 29680 -2410
rect 29770 -2650 30010 -2410
rect 30100 -2650 30340 -2410
rect 30430 -2650 30670 -2410
rect 30760 -2650 31000 -2410
rect 31090 -2650 31330 -2410
rect 31420 -2650 31660 -2410
rect 31750 -2650 31990 -2410
rect 32080 -2650 32320 -2410
rect 32410 -2650 32650 -2410
rect 32740 -2650 32980 -2410
rect 33070 -2650 33310 -2410
rect 33400 -2650 33640 -2410
rect 33730 -2650 33970 -2410
rect 34060 -2650 34300 -2410
rect 34390 -2650 34630 -2410
rect 34720 -2650 34960 -2410
rect 35050 -2650 35290 -2410
rect 28780 -2980 29020 -2740
rect 29110 -2980 29350 -2740
rect 29440 -2980 29680 -2740
rect 29770 -2980 30010 -2740
rect 30100 -2980 30340 -2740
rect 30430 -2980 30670 -2740
rect 30760 -2980 31000 -2740
rect 31090 -2980 31330 -2740
rect 31420 -2980 31660 -2740
rect 31750 -2980 31990 -2740
rect 32080 -2980 32320 -2740
rect 32410 -2980 32650 -2740
rect 32740 -2980 32980 -2740
rect 33070 -2980 33310 -2740
rect 33400 -2980 33640 -2740
rect 33730 -2980 33970 -2740
rect 34060 -2980 34300 -2740
rect 34390 -2980 34630 -2740
rect 34720 -2980 34960 -2740
rect 35050 -2980 35290 -2740
rect 28780 -3310 29020 -3070
rect 29110 -3310 29350 -3070
rect 29440 -3310 29680 -3070
rect 29770 -3310 30010 -3070
rect 30100 -3310 30340 -3070
rect 30430 -3310 30670 -3070
rect 30760 -3310 31000 -3070
rect 31090 -3310 31330 -3070
rect 31420 -3310 31660 -3070
rect 31750 -3310 31990 -3070
rect 32080 -3310 32320 -3070
rect 32410 -3310 32650 -3070
rect 32740 -3310 32980 -3070
rect 33070 -3310 33310 -3070
rect 33400 -3310 33640 -3070
rect 33730 -3310 33970 -3070
rect 34060 -3310 34300 -3070
rect 34390 -3310 34630 -3070
rect 34720 -3310 34960 -3070
rect 35050 -3310 35290 -3070
rect 28780 -3640 29020 -3400
rect 29110 -3640 29350 -3400
rect 29440 -3640 29680 -3400
rect 29770 -3640 30010 -3400
rect 30100 -3640 30340 -3400
rect 30430 -3640 30670 -3400
rect 30760 -3640 31000 -3400
rect 31090 -3640 31330 -3400
rect 31420 -3640 31660 -3400
rect 31750 -3640 31990 -3400
rect 32080 -3640 32320 -3400
rect 32410 -3640 32650 -3400
rect 32740 -3640 32980 -3400
rect 33070 -3640 33310 -3400
rect 33400 -3640 33640 -3400
rect 33730 -3640 33970 -3400
rect 34060 -3640 34300 -3400
rect 34390 -3640 34630 -3400
rect 34720 -3640 34960 -3400
rect 35050 -3640 35290 -3400
rect 28780 -3970 29020 -3730
rect 29110 -3970 29350 -3730
rect 29440 -3970 29680 -3730
rect 29770 -3970 30010 -3730
rect 30100 -3970 30340 -3730
rect 30430 -3970 30670 -3730
rect 30760 -3970 31000 -3730
rect 31090 -3970 31330 -3730
rect 31420 -3970 31660 -3730
rect 31750 -3970 31990 -3730
rect 32080 -3970 32320 -3730
rect 32410 -3970 32650 -3730
rect 32740 -3970 32980 -3730
rect 33070 -3970 33310 -3730
rect 33400 -3970 33640 -3730
rect 33730 -3970 33970 -3730
rect 34060 -3970 34300 -3730
rect 34390 -3970 34630 -3730
rect 34720 -3970 34960 -3730
rect 35050 -3970 35290 -3730
rect -1650 -4500 -1410 -4260
rect -1320 -4500 -1080 -4260
rect -990 -4500 -750 -4260
rect -660 -4500 -420 -4260
rect -1650 -4830 -1410 -4590
rect -1320 -4830 -1080 -4590
rect -990 -4830 -750 -4590
rect -660 -4830 -420 -4590
rect -1650 -5160 -1410 -4920
rect -1320 -5160 -1080 -4920
rect -990 -5160 -750 -4920
rect -660 -5160 -420 -4920
rect -1650 -5490 -1410 -5250
rect -1320 -5490 -1080 -5250
rect -990 -5490 -750 -5250
rect -660 -5490 -420 -5250
rect 28780 -4300 29020 -4060
rect 29110 -4300 29350 -4060
rect 29440 -4300 29680 -4060
rect 29770 -4300 30010 -4060
rect 30100 -4300 30340 -4060
rect 30430 -4300 30670 -4060
rect 30760 -4300 31000 -4060
rect 31090 -4300 31330 -4060
rect 31420 -4300 31660 -4060
rect 31750 -4300 31990 -4060
rect 32080 -4300 32320 -4060
rect 32410 -4300 32650 -4060
rect 32740 -4300 32980 -4060
rect 33070 -4300 33310 -4060
rect 33400 -4300 33640 -4060
rect 33730 -4300 33970 -4060
rect 34060 -4300 34300 -4060
rect 34390 -4300 34630 -4060
rect 34720 -4300 34960 -4060
rect 35050 -4300 35290 -4060
rect 28780 -4630 29020 -4390
rect 29110 -4630 29350 -4390
rect 29440 -4630 29680 -4390
rect 29770 -4630 30010 -4390
rect 30100 -4630 30340 -4390
rect 30430 -4630 30670 -4390
rect 30760 -4630 31000 -4390
rect 31090 -4630 31330 -4390
rect 31420 -4630 31660 -4390
rect 31750 -4630 31990 -4390
rect 32080 -4630 32320 -4390
rect 32410 -4630 32650 -4390
rect 32740 -4630 32980 -4390
rect 33070 -4630 33310 -4390
rect 33400 -4630 33640 -4390
rect 33730 -4630 33970 -4390
rect 34060 -4630 34300 -4390
rect 34390 -4630 34630 -4390
rect 34720 -4630 34960 -4390
rect 35050 -4630 35290 -4390
rect 28780 -4960 29020 -4720
rect 29110 -4960 29350 -4720
rect 29440 -4960 29680 -4720
rect 29770 -4960 30010 -4720
rect 30100 -4960 30340 -4720
rect 30430 -4960 30670 -4720
rect 30760 -4960 31000 -4720
rect 31090 -4960 31330 -4720
rect 31420 -4960 31660 -4720
rect 31750 -4960 31990 -4720
rect 32080 -4960 32320 -4720
rect 32410 -4960 32650 -4720
rect 32740 -4960 32980 -4720
rect 33070 -4960 33310 -4720
rect 33400 -4960 33640 -4720
rect 33730 -4960 33970 -4720
rect 34060 -4960 34300 -4720
rect 34390 -4960 34630 -4720
rect 34720 -4960 34960 -4720
rect 35050 -4960 35290 -4720
rect 28780 -5290 29020 -5050
rect 29110 -5290 29350 -5050
rect 29440 -5290 29680 -5050
rect 29770 -5290 30010 -5050
rect 30100 -5290 30340 -5050
rect 30430 -5290 30670 -5050
rect 30760 -5290 31000 -5050
rect 31090 -5290 31330 -5050
rect 31420 -5290 31660 -5050
rect 31750 -5290 31990 -5050
rect 32080 -5290 32320 -5050
rect 32410 -5290 32650 -5050
rect 32740 -5290 32980 -5050
rect 33070 -5290 33310 -5050
rect 33400 -5290 33640 -5050
rect 33730 -5290 33970 -5050
rect 34060 -5290 34300 -5050
rect 34390 -5290 34630 -5050
rect 34720 -5290 34960 -5050
rect 35050 -5290 35290 -5050
rect 28780 -5620 29020 -5380
rect 29110 -5620 29350 -5380
rect 29440 -5620 29680 -5380
rect 29770 -5620 30010 -5380
rect 30100 -5620 30340 -5380
rect 30430 -5620 30670 -5380
rect 30760 -5620 31000 -5380
rect 31090 -5620 31330 -5380
rect 31420 -5620 31660 -5380
rect 31750 -5620 31990 -5380
rect 32080 -5620 32320 -5380
rect 32410 -5620 32650 -5380
rect 32740 -5620 32980 -5380
rect 33070 -5620 33310 -5380
rect 33400 -5620 33640 -5380
rect 33730 -5620 33970 -5380
rect 34060 -5620 34300 -5380
rect 34390 -5620 34630 -5380
rect 34720 -5620 34960 -5380
rect 35050 -5620 35290 -5380
rect 28780 -5950 29020 -5710
rect 29110 -5950 29350 -5710
rect 29440 -5950 29680 -5710
rect 29770 -5950 30010 -5710
rect 30100 -5950 30340 -5710
rect 30430 -5950 30670 -5710
rect 30760 -5950 31000 -5710
rect 31090 -5950 31330 -5710
rect 31420 -5950 31660 -5710
rect 31750 -5950 31990 -5710
rect 32080 -5950 32320 -5710
rect 32410 -5950 32650 -5710
rect 32740 -5950 32980 -5710
rect 33070 -5950 33310 -5710
rect 33400 -5950 33640 -5710
rect 33730 -5950 33970 -5710
rect 34060 -5950 34300 -5710
rect 34390 -5950 34630 -5710
rect 34720 -5950 34960 -5710
rect 35050 -5950 35290 -5710
rect 28780 -6280 29020 -6040
rect 29110 -6280 29350 -6040
rect 29440 -6280 29680 -6040
rect 29770 -6280 30010 -6040
rect 30100 -6280 30340 -6040
rect 30430 -6280 30670 -6040
rect 30760 -6280 31000 -6040
rect 31090 -6280 31330 -6040
rect 31420 -6280 31660 -6040
rect 31750 -6280 31990 -6040
rect 32080 -6280 32320 -6040
rect 32410 -6280 32650 -6040
rect 32740 -6280 32980 -6040
rect 33070 -6280 33310 -6040
rect 33400 -6280 33640 -6040
rect 33730 -6280 33970 -6040
rect 34060 -6280 34300 -6040
rect 34390 -6280 34630 -6040
rect 34720 -6280 34960 -6040
rect 35050 -6280 35290 -6040
rect -1650 -7900 -1410 -7660
rect -1320 -7900 -1080 -7660
rect -990 -7900 -750 -7660
rect -660 -7900 -420 -7660
rect -1650 -8230 -1410 -7990
rect -1320 -8230 -1080 -7990
rect -990 -8230 -750 -7990
rect -660 -8230 -420 -7990
rect -1650 -8560 -1410 -8320
rect -1320 -8560 -1080 -8320
rect -990 -8560 -750 -8320
rect -660 -8560 -420 -8320
rect -1650 -8890 -1410 -8650
rect -1320 -8890 -1080 -8650
rect -990 -8890 -750 -8650
rect -660 -8890 -420 -8650
<< metal4 >>
rect 7020 21140 7290 21300
rect -5020 20790 7290 21140
rect -5020 20550 -4670 20790
rect -4430 20550 -4340 20790
rect -4100 20550 -4010 20790
rect -3770 20550 -3680 20790
rect -3440 20550 -3350 20790
rect -3110 20550 -3020 20790
rect -2780 20550 -2690 20790
rect -2450 20550 -2360 20790
rect -2120 20550 -2030 20790
rect -1790 20550 -1700 20790
rect -1460 20550 -1370 20790
rect -1130 20550 -1040 20790
rect -800 20550 -710 20790
rect -470 20550 -380 20790
rect -140 20550 -50 20790
rect 190 20550 280 20790
rect 520 20550 610 20790
rect 850 20550 940 20790
rect 1180 20550 1270 20790
rect 1510 20550 1600 20790
rect 1840 20550 1930 20790
rect 2170 20550 2260 20790
rect 2500 20550 2590 20790
rect 2830 20550 2920 20790
rect 3160 20550 3250 20790
rect 3490 20550 3580 20790
rect 3820 20550 3910 20790
rect 4150 20550 4240 20790
rect 4480 20550 4570 20790
rect 4810 20550 4900 20790
rect 5140 20550 5230 20790
rect 5470 20550 5560 20790
rect 5800 20550 5890 20790
rect 6130 20550 6220 20790
rect 6460 20550 6550 20790
rect 6790 20550 6880 20790
rect 7120 20550 7290 20790
rect -5020 20460 7290 20550
rect -5020 20220 -4670 20460
rect -4430 20220 -4340 20460
rect -4100 20220 -4010 20460
rect -3770 20220 -3680 20460
rect -3440 20220 -3350 20460
rect -3110 20220 -3020 20460
rect -2780 20220 -2690 20460
rect -2450 20220 -2360 20460
rect -2120 20220 -2030 20460
rect -1790 20220 -1700 20460
rect -1460 20220 -1370 20460
rect -1130 20220 -1040 20460
rect -800 20220 -710 20460
rect -470 20220 -380 20460
rect -140 20220 -50 20460
rect 190 20220 280 20460
rect 520 20220 610 20460
rect 850 20220 940 20460
rect 1180 20220 1270 20460
rect 1510 20220 1600 20460
rect 1840 20220 1930 20460
rect 2170 20220 2260 20460
rect 2500 20220 2590 20460
rect 2830 20220 2920 20460
rect 3160 20220 3250 20460
rect 3490 20220 3580 20460
rect 3820 20220 3910 20460
rect 4150 20220 4240 20460
rect 4480 20220 4570 20460
rect 4810 20220 4900 20460
rect 5140 20220 5230 20460
rect 5470 20220 5560 20460
rect 5800 20220 5890 20460
rect 6130 20220 6220 20460
rect 6460 20220 6550 20460
rect 6790 20220 6880 20460
rect 7120 20220 7290 20460
rect -5020 20130 7290 20220
rect -5020 19890 -4670 20130
rect -4430 19890 -4340 20130
rect -4100 19890 -4010 20130
rect -3770 19890 -3680 20130
rect -3440 19890 -3350 20130
rect -3110 19890 -3020 20130
rect -2780 19890 -2690 20130
rect -2450 19890 -2360 20130
rect -2120 19890 -2030 20130
rect -1790 19890 -1700 20130
rect -1460 19890 -1370 20130
rect -1130 19890 -1040 20130
rect -800 19890 -710 20130
rect -470 19890 -380 20130
rect -140 19890 -50 20130
rect 190 19890 280 20130
rect 520 19890 610 20130
rect 850 19890 940 20130
rect 1180 19890 1270 20130
rect 1510 19890 1600 20130
rect 1840 19890 1930 20130
rect 2170 19890 2260 20130
rect 2500 19890 2590 20130
rect 2830 19890 2920 20130
rect 3160 19890 3250 20130
rect 3490 19890 3580 20130
rect 3820 19890 3910 20130
rect 4150 19890 4240 20130
rect 4480 19890 4570 20130
rect 4810 19890 4900 20130
rect 5140 19890 5230 20130
rect 5470 19890 5560 20130
rect 5800 19890 5890 20130
rect 6130 19890 6220 20130
rect 6460 19890 6550 20130
rect 6790 19890 6880 20130
rect 7120 19890 7290 20130
rect -5020 19800 7290 19890
rect -5020 19560 -4670 19800
rect -4430 19560 -4340 19800
rect -4100 19560 -4010 19800
rect -3770 19560 -3680 19800
rect -3440 19560 -3350 19800
rect -3110 19560 -3020 19800
rect -2780 19560 -2690 19800
rect -2450 19560 -2360 19800
rect -2120 19560 -2030 19800
rect -1790 19560 -1700 19800
rect -1460 19560 -1370 19800
rect -1130 19560 -1040 19800
rect -800 19560 -710 19800
rect -470 19560 -380 19800
rect -140 19560 -50 19800
rect 190 19560 280 19800
rect 520 19560 610 19800
rect 850 19560 940 19800
rect 1180 19560 1270 19800
rect 1510 19560 1600 19800
rect 1840 19560 1930 19800
rect 2170 19560 2260 19800
rect 2500 19560 2590 19800
rect 2830 19560 2920 19800
rect 3160 19560 3250 19800
rect 3490 19560 3580 19800
rect 3820 19560 3910 19800
rect 4150 19560 4240 19800
rect 4480 19560 4570 19800
rect 4810 19560 4900 19800
rect 5140 19560 5230 19800
rect 5470 19560 5560 19800
rect 5800 19560 5890 19800
rect 6130 19560 6220 19800
rect 6460 19560 6550 19800
rect 6790 19560 6880 19800
rect 7120 19560 7290 19800
rect -5020 19470 7290 19560
rect -5020 19230 -4670 19470
rect -4430 19230 -4340 19470
rect -4100 19230 -4010 19470
rect -3770 19230 -3680 19470
rect -3440 19230 -3350 19470
rect -3110 19230 -3020 19470
rect -2780 19230 -2690 19470
rect -2450 19230 -2360 19470
rect -2120 19230 -2030 19470
rect -1790 19230 -1700 19470
rect -1460 19230 -1370 19470
rect -1130 19230 -1040 19470
rect -800 19230 -710 19470
rect -470 19230 -380 19470
rect -140 19230 -50 19470
rect 190 19230 280 19470
rect 520 19230 610 19470
rect 850 19230 940 19470
rect 1180 19230 1270 19470
rect 1510 19230 1600 19470
rect 1840 19230 1930 19470
rect 2170 19230 2260 19470
rect 2500 19230 2590 19470
rect 2830 19230 2920 19470
rect 3160 19230 3250 19470
rect 3490 19230 3580 19470
rect 3820 19230 3910 19470
rect 4150 19230 4240 19470
rect 4480 19230 4570 19470
rect 4810 19230 4900 19470
rect 5140 19230 5230 19470
rect 5470 19230 5560 19470
rect 5800 19230 5890 19470
rect 6130 19230 6220 19470
rect 6460 19230 6550 19470
rect 6790 19230 6880 19470
rect 7120 19230 7290 19470
rect -5020 19140 7290 19230
rect -5020 18900 -4670 19140
rect -4430 18900 -4340 19140
rect -4100 18900 -4010 19140
rect -3770 18900 -3680 19140
rect -3440 18900 -3350 19140
rect -3110 18900 -3020 19140
rect -2780 18900 -2690 19140
rect -2450 18900 -2360 19140
rect -2120 18900 -2030 19140
rect -1790 18900 -1700 19140
rect -1460 18900 -1370 19140
rect -1130 18900 -1040 19140
rect -800 18900 -710 19140
rect -470 18900 -380 19140
rect -140 18900 -50 19140
rect 190 18900 280 19140
rect 520 18900 610 19140
rect 850 18900 940 19140
rect 1180 18900 1270 19140
rect 1510 18900 1600 19140
rect 1840 18900 1930 19140
rect 2170 18900 2260 19140
rect 2500 18900 2590 19140
rect 2830 18900 2920 19140
rect 3160 18900 3250 19140
rect 3490 18900 3580 19140
rect 3820 18900 3910 19140
rect 4150 18900 4240 19140
rect 4480 18900 4570 19140
rect 4810 18900 4900 19140
rect 5140 18900 5230 19140
rect 5470 18900 5560 19140
rect 5800 18900 5890 19140
rect 6130 18900 6220 19140
rect 6460 18900 6550 19140
rect 6790 18900 6880 19140
rect 7120 18900 7290 19140
rect -5020 18810 7290 18900
rect -5020 18570 -4670 18810
rect -4430 18570 -4340 18810
rect -4100 18570 -4010 18810
rect -3770 18570 -3680 18810
rect -3440 18570 -3350 18810
rect -3110 18570 -3020 18810
rect -2780 18570 -2690 18810
rect -2450 18570 -2360 18810
rect -2120 18570 -2030 18810
rect -1790 18570 -1700 18810
rect -1460 18570 -1370 18810
rect -1130 18570 -1040 18810
rect -800 18570 -710 18810
rect -470 18570 -380 18810
rect -140 18570 -50 18810
rect 190 18570 280 18810
rect 520 18570 610 18810
rect 850 18570 940 18810
rect 1180 18570 1270 18810
rect 1510 18570 1600 18810
rect 1840 18570 1930 18810
rect 2170 18570 2260 18810
rect 2500 18570 2590 18810
rect 2830 18570 2920 18810
rect 3160 18570 3250 18810
rect 3490 18570 3580 18810
rect 3820 18570 3910 18810
rect 4150 18570 4240 18810
rect 4480 18570 4570 18810
rect 4810 18570 4900 18810
rect 5140 18570 5230 18810
rect 5470 18570 5560 18810
rect 5800 18570 5890 18810
rect 6130 18570 6220 18810
rect 6460 18570 6550 18810
rect 6790 18570 6880 18810
rect 7120 18570 7290 18810
rect -5020 18480 7290 18570
rect -5020 18240 -4670 18480
rect -4430 18240 -4340 18480
rect -4100 18240 -4010 18480
rect -3770 18240 -3680 18480
rect -3440 18240 -3350 18480
rect -3110 18240 -3020 18480
rect -2780 18240 -2690 18480
rect -2450 18240 -2360 18480
rect -2120 18240 -2030 18480
rect -1790 18240 -1700 18480
rect -1460 18240 -1370 18480
rect -1130 18240 -1040 18480
rect -800 18240 -710 18480
rect -470 18240 -380 18480
rect -140 18240 -50 18480
rect 190 18240 280 18480
rect 520 18240 610 18480
rect 850 18240 940 18480
rect 1180 18240 1270 18480
rect 1510 18240 1600 18480
rect 1840 18240 1930 18480
rect 2170 18240 2260 18480
rect 2500 18240 2590 18480
rect 2830 18240 2920 18480
rect 3160 18240 3250 18480
rect 3490 18240 3580 18480
rect 3820 18240 3910 18480
rect 4150 18240 4240 18480
rect 4480 18240 4570 18480
rect 4810 18240 4900 18480
rect 5140 18240 5230 18480
rect 5470 18240 5560 18480
rect 5800 18240 5890 18480
rect 6130 18240 6220 18480
rect 6460 18240 6550 18480
rect 6790 18240 6880 18480
rect 7120 18240 7290 18480
rect -5020 18150 7290 18240
rect -5020 17910 -4670 18150
rect -4430 17910 -4340 18150
rect -4100 17910 -4010 18150
rect -3770 17910 -3680 18150
rect -3440 17910 -3350 18150
rect -3110 17910 -3020 18150
rect -2780 17910 -2690 18150
rect -2450 17910 -2360 18150
rect -2120 17910 -2030 18150
rect -1790 17910 -1700 18150
rect -1460 17910 -1370 18150
rect -1130 17910 -1040 18150
rect -800 17910 -710 18150
rect -470 17910 -380 18150
rect -140 17910 -50 18150
rect 190 17910 280 18150
rect 520 17910 610 18150
rect 850 17910 940 18150
rect 1180 17910 1270 18150
rect 1510 17910 1600 18150
rect 1840 17910 1930 18150
rect 2170 17910 2260 18150
rect 2500 17910 2590 18150
rect 2830 17910 2920 18150
rect 3160 17910 3250 18150
rect 3490 17910 3580 18150
rect 3820 17910 3910 18150
rect 4150 17910 4240 18150
rect 4480 17910 4570 18150
rect 4810 17910 4900 18150
rect 5140 17910 5230 18150
rect 5470 17910 5560 18150
rect 5800 17910 5890 18150
rect 6130 17910 6220 18150
rect 6460 17910 6550 18150
rect 6790 17910 6880 18150
rect 7120 17910 7290 18150
rect -5020 17820 7290 17910
rect -5020 17580 -4670 17820
rect -4430 17580 -4340 17820
rect -4100 17580 -4010 17820
rect -3770 17580 -3680 17820
rect -3440 17580 -3350 17820
rect -3110 17580 -3020 17820
rect -2780 17580 -2690 17820
rect -2450 17580 -2360 17820
rect -2120 17580 -2030 17820
rect -1790 17580 -1700 17820
rect -1460 17580 -1370 17820
rect -1130 17580 -1040 17820
rect -800 17580 -710 17820
rect -470 17580 -380 17820
rect -140 17580 -50 17820
rect 190 17580 280 17820
rect 520 17580 610 17820
rect 850 17580 940 17820
rect 1180 17580 1270 17820
rect 1510 17580 1600 17820
rect 1840 17580 1930 17820
rect 2170 17580 2260 17820
rect 2500 17580 2590 17820
rect 2830 17580 2920 17820
rect 3160 17580 3250 17820
rect 3490 17580 3580 17820
rect 3820 17580 3910 17820
rect 4150 17580 4240 17820
rect 4480 17580 4570 17820
rect 4810 17580 4900 17820
rect 5140 17580 5230 17820
rect 5470 17580 5560 17820
rect 5800 17580 5890 17820
rect 6130 17580 6220 17820
rect 6460 17580 6550 17820
rect 6790 17580 6880 17820
rect 7120 17580 7290 17820
rect -5020 17490 7290 17580
rect -5020 17250 -4670 17490
rect -4430 17250 -4340 17490
rect -4100 17250 -4010 17490
rect -3770 17250 -3680 17490
rect -3440 17250 -3350 17490
rect -3110 17250 -3020 17490
rect -2780 17250 -2690 17490
rect -2450 17250 -2360 17490
rect -2120 17250 -2030 17490
rect -1790 17250 -1700 17490
rect -1460 17250 -1370 17490
rect -1130 17250 -1040 17490
rect -800 17250 -710 17490
rect -470 17250 -380 17490
rect -140 17250 -50 17490
rect 190 17250 280 17490
rect 520 17250 610 17490
rect 850 17250 940 17490
rect 1180 17250 1270 17490
rect 1510 17250 1600 17490
rect 1840 17250 1930 17490
rect 2170 17250 2260 17490
rect 2500 17250 2590 17490
rect 2830 17250 2920 17490
rect 3160 17250 3250 17490
rect 3490 17250 3580 17490
rect 3820 17250 3910 17490
rect 4150 17250 4240 17490
rect 4480 17250 4570 17490
rect 4810 17250 4900 17490
rect 5140 17250 5230 17490
rect 5470 17250 5560 17490
rect 5800 17250 5890 17490
rect 6130 17250 6220 17490
rect 6460 17250 6550 17490
rect 6790 17250 6880 17490
rect 7120 17250 7290 17490
rect -5020 17160 7290 17250
rect -5020 16920 -4670 17160
rect -4430 16920 -4340 17160
rect -4100 16920 -4010 17160
rect -3770 16920 -3680 17160
rect -3440 16920 -3350 17160
rect -3110 16920 -3020 17160
rect -2780 16920 -2690 17160
rect -2450 16920 -2360 17160
rect -2120 16920 -2030 17160
rect -1790 16920 -1700 17160
rect -1460 16920 -1370 17160
rect -1130 16920 -1040 17160
rect -800 16920 -710 17160
rect -470 16920 -380 17160
rect -140 16920 -50 17160
rect 190 16920 280 17160
rect 520 16920 610 17160
rect 850 16920 940 17160
rect 1180 16920 1270 17160
rect 1510 16920 1600 17160
rect 1840 16920 1930 17160
rect 2170 16920 2260 17160
rect 2500 16920 2590 17160
rect 2830 16920 2920 17160
rect 3160 16920 3250 17160
rect 3490 16920 3580 17160
rect 3820 16920 3910 17160
rect 4150 16920 4240 17160
rect 4480 16920 4570 17160
rect 4810 16920 4900 17160
rect 5140 16920 5230 17160
rect 5470 16920 5560 17160
rect 5800 16920 5890 17160
rect 6130 16920 6220 17160
rect 6460 16920 6550 17160
rect 6790 16920 6880 17160
rect 7120 16920 7290 17160
rect -5020 16830 7290 16920
rect -5020 16590 -4670 16830
rect -4430 16590 -4340 16830
rect -4100 16590 -4010 16830
rect -3770 16590 -3680 16830
rect -3440 16590 -3350 16830
rect -3110 16590 -3020 16830
rect -2780 16590 -2690 16830
rect -2450 16590 -2360 16830
rect -2120 16590 -2030 16830
rect -1790 16590 -1700 16830
rect -1460 16590 -1370 16830
rect -1130 16590 -1040 16830
rect -800 16590 -710 16830
rect -470 16590 -380 16830
rect -140 16590 -50 16830
rect 190 16590 280 16830
rect 520 16590 610 16830
rect 850 16590 940 16830
rect 1180 16590 1270 16830
rect 1510 16590 1600 16830
rect 1840 16590 1930 16830
rect 2170 16590 2260 16830
rect 2500 16590 2590 16830
rect 2830 16590 2920 16830
rect 3160 16590 3250 16830
rect 3490 16590 3580 16830
rect 3820 16590 3910 16830
rect 4150 16590 4240 16830
rect 4480 16590 4570 16830
rect 4810 16590 4900 16830
rect 5140 16590 5230 16830
rect 5470 16590 5560 16830
rect 5800 16590 5890 16830
rect 6130 16590 6220 16830
rect 6460 16590 6550 16830
rect 6790 16590 6880 16830
rect 7120 16590 7290 16830
rect -5020 16500 7290 16590
rect -5020 16260 -4670 16500
rect -4430 16260 -4340 16500
rect -4100 16260 -4010 16500
rect -3770 16260 -3680 16500
rect -3440 16260 -3350 16500
rect -3110 16260 -3020 16500
rect -2780 16260 -2690 16500
rect -2450 16260 -2360 16500
rect -2120 16260 -2030 16500
rect -1790 16260 -1700 16500
rect -1460 16260 -1370 16500
rect -1130 16260 -1040 16500
rect -800 16260 -710 16500
rect -470 16260 -380 16500
rect -140 16260 -50 16500
rect 190 16260 280 16500
rect 520 16260 610 16500
rect 850 16260 940 16500
rect 1180 16260 1270 16500
rect 1510 16260 1600 16500
rect 1840 16260 1930 16500
rect 2170 16260 2260 16500
rect 2500 16260 2590 16500
rect 2830 16260 2920 16500
rect 3160 16260 3250 16500
rect 3490 16260 3580 16500
rect 3820 16260 3910 16500
rect 4150 16260 4240 16500
rect 4480 16260 4570 16500
rect 4810 16260 4900 16500
rect 5140 16260 5230 16500
rect 5470 16260 5560 16500
rect 5800 16260 5890 16500
rect 6130 16260 6220 16500
rect 6460 16260 6550 16500
rect 6790 16260 6880 16500
rect 7120 16260 7290 16500
rect -5020 16170 7290 16260
rect -5020 15930 -4670 16170
rect -4430 15930 -4340 16170
rect -4100 15930 -4010 16170
rect -3770 15930 -3680 16170
rect -3440 15930 -3350 16170
rect -3110 15930 -3020 16170
rect -2780 15930 -2690 16170
rect -2450 15930 -2360 16170
rect -2120 15930 -2030 16170
rect -1790 15930 -1700 16170
rect -1460 15930 -1370 16170
rect -1130 15930 -1040 16170
rect -800 15930 -710 16170
rect -470 15930 -380 16170
rect -140 15930 -50 16170
rect 190 15930 280 16170
rect 520 15930 610 16170
rect 850 15930 940 16170
rect 1180 15930 1270 16170
rect 1510 15930 1600 16170
rect 1840 15930 1930 16170
rect 2170 15930 2260 16170
rect 2500 15930 2590 16170
rect 2830 15930 2920 16170
rect 3160 15930 3250 16170
rect 3490 15930 3580 16170
rect 3820 15930 3910 16170
rect 4150 15930 4240 16170
rect 4480 15930 4570 16170
rect 4810 15930 4900 16170
rect 5140 15930 5230 16170
rect 5470 15930 5560 16170
rect 5800 15930 5890 16170
rect 6130 15930 6220 16170
rect 6460 15930 6550 16170
rect 6790 15930 6880 16170
rect 7120 15930 7290 16170
rect -5020 15840 7290 15930
rect -5020 15600 -4670 15840
rect -4430 15600 -4340 15840
rect -4100 15600 -4010 15840
rect -3770 15600 -3680 15840
rect -3440 15600 -3350 15840
rect -3110 15600 -3020 15840
rect -2780 15600 -2690 15840
rect -2450 15600 -2360 15840
rect -2120 15600 -2030 15840
rect -1790 15600 -1700 15840
rect -1460 15600 -1370 15840
rect -1130 15600 -1040 15840
rect -800 15600 -710 15840
rect -470 15600 -380 15840
rect -140 15600 -50 15840
rect 190 15600 280 15840
rect 520 15600 610 15840
rect 850 15600 940 15840
rect 1180 15600 1270 15840
rect 1510 15600 1600 15840
rect 1840 15600 1930 15840
rect 2170 15600 2260 15840
rect 2500 15600 2590 15840
rect 2830 15600 2920 15840
rect 3160 15600 3250 15840
rect 3490 15600 3580 15840
rect 3820 15600 3910 15840
rect 4150 15600 4240 15840
rect 4480 15600 4570 15840
rect 4810 15600 4900 15840
rect 5140 15600 5230 15840
rect 5470 15600 5560 15840
rect 5800 15600 5890 15840
rect 6130 15600 6220 15840
rect 6460 15600 6550 15840
rect 6790 15600 6880 15840
rect 7120 15600 7290 15840
rect -5020 15510 7290 15600
rect -5020 15270 -4670 15510
rect -4430 15270 -4340 15510
rect -4100 15270 -4010 15510
rect -3770 15270 -3680 15510
rect -3440 15270 -3350 15510
rect -3110 15270 -3020 15510
rect -2780 15270 -2690 15510
rect -2450 15270 -2360 15510
rect -2120 15270 -2030 15510
rect -1790 15270 -1700 15510
rect -1460 15270 -1370 15510
rect -1130 15270 -1040 15510
rect -800 15270 -710 15510
rect -470 15270 -380 15510
rect -140 15270 -50 15510
rect 190 15270 280 15510
rect 520 15270 610 15510
rect 850 15270 940 15510
rect 1180 15270 1270 15510
rect 1510 15270 1600 15510
rect 1840 15270 1930 15510
rect 2170 15270 2260 15510
rect 2500 15270 2590 15510
rect 2830 15270 2920 15510
rect 3160 15270 3250 15510
rect 3490 15270 3580 15510
rect 3820 15270 3910 15510
rect 4150 15270 4240 15510
rect 4480 15270 4570 15510
rect 4810 15270 4900 15510
rect 5140 15270 5230 15510
rect 5470 15270 5560 15510
rect 5800 15270 5890 15510
rect 6130 15270 6220 15510
rect 6460 15270 6550 15510
rect 6790 15270 6880 15510
rect 7120 15270 7290 15510
rect -5020 15180 7290 15270
rect -5020 14940 -4670 15180
rect -4430 14940 -4340 15180
rect -4100 14940 -4010 15180
rect -3770 14940 -3680 15180
rect -3440 14940 -3350 15180
rect -3110 14940 -3020 15180
rect -2780 14940 -2690 15180
rect -2450 14940 -2360 15180
rect -2120 14940 -2030 15180
rect -1790 14940 -1700 15180
rect -1460 14940 -1370 15180
rect -1130 14940 -1040 15180
rect -800 14940 -710 15180
rect -470 14940 -380 15180
rect -140 14940 -50 15180
rect 190 14940 280 15180
rect 520 14940 610 15180
rect 850 14940 940 15180
rect 1180 14940 1270 15180
rect 1510 14940 1600 15180
rect 1840 14940 1930 15180
rect 2170 14940 2260 15180
rect 2500 14940 2590 15180
rect 2830 14940 2920 15180
rect 3160 14940 3250 15180
rect 3490 14940 3580 15180
rect 3820 14940 3910 15180
rect 4150 14940 4240 15180
rect 4480 14940 4570 15180
rect 4810 14940 4900 15180
rect 5140 14940 5230 15180
rect 5470 14940 5560 15180
rect 5800 14940 5890 15180
rect 6130 14940 6220 15180
rect 6460 14940 6550 15180
rect 6790 14940 6880 15180
rect 7120 14940 7290 15180
rect -5020 14850 7290 14940
rect -5020 14610 -4670 14850
rect -4430 14610 -4340 14850
rect -4100 14610 -4010 14850
rect -3770 14610 -3680 14850
rect -3440 14610 -3350 14850
rect -3110 14610 -3020 14850
rect -2780 14610 -2690 14850
rect -2450 14610 -2360 14850
rect -2120 14610 -2030 14850
rect -1790 14610 -1700 14850
rect -1460 14610 -1370 14850
rect -1130 14610 -1040 14850
rect -800 14610 -710 14850
rect -470 14610 -380 14850
rect -140 14610 -50 14850
rect 190 14610 280 14850
rect 520 14610 610 14850
rect 850 14610 940 14850
rect 1180 14610 1270 14850
rect 1510 14610 1600 14850
rect 1840 14610 1930 14850
rect 2170 14610 2260 14850
rect 2500 14610 2590 14850
rect 2830 14610 2920 14850
rect 3160 14610 3250 14850
rect 3490 14610 3580 14850
rect 3820 14610 3910 14850
rect 4150 14610 4240 14850
rect 4480 14610 4570 14850
rect 4810 14610 4900 14850
rect 5140 14610 5230 14850
rect 5470 14610 5560 14850
rect 5800 14610 5890 14850
rect 6130 14610 6220 14850
rect 6460 14610 6550 14850
rect 6790 14610 6880 14850
rect 7120 14610 7290 14850
rect -5020 14520 7290 14610
rect -5020 14280 -4670 14520
rect -4430 14280 -4340 14520
rect -4100 14280 -4010 14520
rect -3770 14280 -3680 14520
rect -3440 14280 -3350 14520
rect -3110 14280 -3020 14520
rect -2780 14280 -2690 14520
rect -2450 14280 -2360 14520
rect -2120 14280 -2030 14520
rect -1790 14280 -1700 14520
rect -1460 14280 -1370 14520
rect -1130 14280 -1040 14520
rect -800 14280 -710 14520
rect -470 14280 -380 14520
rect -140 14280 -50 14520
rect 190 14280 280 14520
rect 520 14280 610 14520
rect 850 14280 940 14520
rect 1180 14280 1270 14520
rect 1510 14280 1600 14520
rect 1840 14280 1930 14520
rect 2170 14280 2260 14520
rect 2500 14280 2590 14520
rect 2830 14280 2920 14520
rect 3160 14280 3250 14520
rect 3490 14280 3580 14520
rect 3820 14280 3910 14520
rect 4150 14280 4240 14520
rect 4480 14280 4570 14520
rect 4810 14280 4900 14520
rect 5140 14280 5230 14520
rect 5470 14280 5560 14520
rect 5800 14280 5890 14520
rect 6130 14280 6220 14520
rect 6460 14280 6550 14520
rect 6790 14280 6880 14520
rect 7120 14280 7290 14520
rect -5020 14190 7290 14280
rect -5020 13950 -4670 14190
rect -4430 13950 -4340 14190
rect -4100 13950 -4010 14190
rect -3770 13950 -3680 14190
rect -3440 13950 -3350 14190
rect -3110 13950 -3020 14190
rect -2780 13950 -2690 14190
rect -2450 13950 -2360 14190
rect -2120 13950 -2030 14190
rect -1790 13950 -1700 14190
rect -1460 13950 -1370 14190
rect -1130 13950 -1040 14190
rect -800 13950 -710 14190
rect -470 13950 -380 14190
rect -140 13950 -50 14190
rect 190 13950 280 14190
rect 520 13950 610 14190
rect 850 13950 940 14190
rect 1180 13950 1270 14190
rect 1510 13950 1600 14190
rect 1840 13950 1930 14190
rect 2170 13950 2260 14190
rect 2500 13950 2590 14190
rect 2830 13950 2920 14190
rect 3160 13950 3250 14190
rect 3490 13950 3580 14190
rect 3820 13950 3910 14190
rect 4150 13950 4240 14190
rect 4480 13950 4570 14190
rect 4810 13950 4900 14190
rect 5140 13950 5230 14190
rect 5470 13950 5560 14190
rect 5800 13950 5890 14190
rect 6130 13950 6220 14190
rect 6460 13950 6550 14190
rect 6790 13950 6880 14190
rect 7120 13950 7290 14190
rect -5020 13860 7290 13950
rect -5020 13620 -4670 13860
rect -4430 13620 -4340 13860
rect -4100 13620 -4010 13860
rect -3770 13620 -3680 13860
rect -3440 13620 -3350 13860
rect -3110 13620 -3020 13860
rect -2780 13620 -2690 13860
rect -2450 13620 -2360 13860
rect -2120 13620 -2030 13860
rect -1790 13620 -1700 13860
rect -1460 13620 -1370 13860
rect -1130 13620 -1040 13860
rect -800 13620 -710 13860
rect -470 13620 -380 13860
rect -140 13620 -50 13860
rect 190 13620 280 13860
rect 520 13620 610 13860
rect 850 13620 940 13860
rect 1180 13620 1270 13860
rect 1510 13620 1600 13860
rect 1840 13620 1930 13860
rect 2170 13620 2260 13860
rect 2500 13620 2590 13860
rect 2830 13620 2920 13860
rect 3160 13620 3250 13860
rect 3490 13620 3580 13860
rect 3820 13620 3910 13860
rect 4150 13620 4240 13860
rect 4480 13620 4570 13860
rect 4810 13620 4900 13860
rect 5140 13620 5230 13860
rect 5470 13620 5560 13860
rect 5800 13620 5890 13860
rect 6130 13620 6220 13860
rect 6460 13620 6550 13860
rect 6790 13620 6880 13860
rect 7120 13620 7290 13860
rect -5020 13530 7290 13620
rect -5020 13290 -4670 13530
rect -4430 13290 -4340 13530
rect -4100 13290 -4010 13530
rect -3770 13290 -3680 13530
rect -3440 13290 -3350 13530
rect -3110 13290 -3020 13530
rect -2780 13290 -2690 13530
rect -2450 13290 -2360 13530
rect -2120 13290 -2030 13530
rect -1790 13290 -1700 13530
rect -1460 13290 -1370 13530
rect -1130 13290 -1040 13530
rect -800 13290 -710 13530
rect -470 13290 -380 13530
rect -140 13290 -50 13530
rect 190 13290 280 13530
rect 520 13290 610 13530
rect 850 13290 940 13530
rect 1180 13290 1270 13530
rect 1510 13290 1600 13530
rect 1840 13290 1930 13530
rect 2170 13290 2260 13530
rect 2500 13290 2590 13530
rect 2830 13290 2920 13530
rect 3160 13290 3250 13530
rect 3490 13290 3580 13530
rect 3820 13290 3910 13530
rect 4150 13290 4240 13530
rect 4480 13290 4570 13530
rect 4810 13290 4900 13530
rect 5140 13290 5230 13530
rect 5470 13290 5560 13530
rect 5800 13290 5890 13530
rect 6130 13290 6220 13530
rect 6460 13290 6550 13530
rect 6790 13290 6880 13530
rect 7120 13290 7290 13530
rect -5020 13200 7290 13290
rect -5020 12960 -4670 13200
rect -4430 12960 -4340 13200
rect -4100 12960 -4010 13200
rect -3770 12960 -3680 13200
rect -3440 12960 -3350 13200
rect -3110 12960 -3020 13200
rect -2780 12960 -2690 13200
rect -2450 12960 -2360 13200
rect -2120 12960 -2030 13200
rect -1790 12960 -1700 13200
rect -1460 12960 -1370 13200
rect -1130 12960 -1040 13200
rect -800 12960 -710 13200
rect -470 12960 -380 13200
rect -140 12960 -50 13200
rect 190 12960 280 13200
rect 520 12960 610 13200
rect 850 12960 940 13200
rect 1180 12960 1270 13200
rect 1510 12960 1600 13200
rect 1840 12960 1930 13200
rect 2170 12960 2260 13200
rect 2500 12960 2590 13200
rect 2830 12960 2920 13200
rect 3160 12960 3250 13200
rect 3490 12960 3580 13200
rect 3820 12960 3910 13200
rect 4150 12960 4240 13200
rect 4480 12960 4570 13200
rect 4810 12960 4900 13200
rect 5140 12960 5230 13200
rect 5470 12960 5560 13200
rect 5800 12960 5890 13200
rect 6130 12960 6220 13200
rect 6460 12960 6550 13200
rect 6790 12960 6880 13200
rect 7120 12960 7290 13200
rect -5020 12870 7290 12960
rect -5020 12630 -4670 12870
rect -4430 12630 -4340 12870
rect -4100 12630 -4010 12870
rect -3770 12630 -3680 12870
rect -3440 12630 -3350 12870
rect -3110 12630 -3020 12870
rect -2780 12630 -2690 12870
rect -2450 12630 -2360 12870
rect -2120 12630 -2030 12870
rect -1790 12630 -1700 12870
rect -1460 12630 -1370 12870
rect -1130 12630 -1040 12870
rect -800 12630 -710 12870
rect -470 12630 -380 12870
rect -140 12630 -50 12870
rect 190 12630 280 12870
rect 520 12630 610 12870
rect 850 12630 940 12870
rect 1180 12630 1270 12870
rect 1510 12630 1600 12870
rect 1840 12630 1930 12870
rect 2170 12630 2260 12870
rect 2500 12630 2590 12870
rect 2830 12630 2920 12870
rect 3160 12630 3250 12870
rect 3490 12630 3580 12870
rect 3820 12630 3910 12870
rect 4150 12630 4240 12870
rect 4480 12630 4570 12870
rect 4810 12630 4900 12870
rect 5140 12630 5230 12870
rect 5470 12630 5560 12870
rect 5800 12630 5890 12870
rect 6130 12630 6220 12870
rect 6460 12630 6550 12870
rect 6790 12630 6880 12870
rect 7120 12630 7290 12870
rect -5020 12540 7290 12630
rect -5020 12300 -4670 12540
rect -4430 12300 -4340 12540
rect -4100 12300 -4010 12540
rect -3770 12300 -3680 12540
rect -3440 12300 -3350 12540
rect -3110 12300 -3020 12540
rect -2780 12300 -2690 12540
rect -2450 12300 -2360 12540
rect -2120 12300 -2030 12540
rect -1790 12300 -1700 12540
rect -1460 12300 -1370 12540
rect -1130 12300 -1040 12540
rect -800 12300 -710 12540
rect -470 12300 -380 12540
rect -140 12300 -50 12540
rect 190 12300 280 12540
rect 520 12300 610 12540
rect 850 12300 940 12540
rect 1180 12300 1270 12540
rect 1510 12300 1600 12540
rect 1840 12300 1930 12540
rect 2170 12300 2260 12540
rect 2500 12300 2590 12540
rect 2830 12300 2920 12540
rect 3160 12300 3250 12540
rect 3490 12300 3580 12540
rect 3820 12300 3910 12540
rect 4150 12300 4240 12540
rect 4480 12300 4570 12540
rect 4810 12300 4900 12540
rect 5140 12300 5230 12540
rect 5470 12300 5560 12540
rect 5800 12300 5890 12540
rect 6130 12300 6220 12540
rect 6460 12300 6550 12540
rect 6790 12300 6880 12540
rect 7120 12300 7290 12540
rect -5020 12210 7290 12300
rect -5020 11970 -4670 12210
rect -4430 11970 -4340 12210
rect -4100 11970 -4010 12210
rect -3770 11970 -3680 12210
rect -3440 11970 -3350 12210
rect -3110 11970 -3020 12210
rect -2780 11970 -2690 12210
rect -2450 11970 -2360 12210
rect -2120 11970 -2030 12210
rect -1790 11970 -1700 12210
rect -1460 11970 -1370 12210
rect -1130 11970 -1040 12210
rect -800 11970 -710 12210
rect -470 11970 -380 12210
rect -140 11970 -50 12210
rect 190 11970 280 12210
rect 520 11970 610 12210
rect 850 11970 940 12210
rect 1180 11970 1270 12210
rect 1510 11970 1600 12210
rect 1840 11970 1930 12210
rect 2170 11970 2260 12210
rect 2500 11970 2590 12210
rect 2830 11970 2920 12210
rect 3160 11970 3250 12210
rect 3490 11970 3580 12210
rect 3820 11970 3910 12210
rect 4150 11970 4240 12210
rect 4480 11970 4570 12210
rect 4810 11970 4900 12210
rect 5140 11970 5230 12210
rect 5470 11970 5560 12210
rect 5800 11970 5890 12210
rect 6130 11970 6220 12210
rect 6460 11970 6550 12210
rect 6790 11970 6880 12210
rect 7120 11970 7290 12210
rect -5020 11880 7290 11970
rect -5020 11640 -4670 11880
rect -4430 11640 -4340 11880
rect -4100 11640 -4010 11880
rect -3770 11640 -3680 11880
rect -3440 11640 -3350 11880
rect -3110 11640 -3020 11880
rect -2780 11640 -2690 11880
rect -2450 11640 -2360 11880
rect -2120 11640 -2030 11880
rect -1790 11640 -1700 11880
rect -1460 11640 -1370 11880
rect -1130 11640 -1040 11880
rect -800 11640 -710 11880
rect -470 11640 -380 11880
rect -140 11640 -50 11880
rect 190 11640 280 11880
rect 520 11640 610 11880
rect 850 11640 940 11880
rect 1180 11640 1270 11880
rect 1510 11640 1600 11880
rect 1840 11640 1930 11880
rect 2170 11640 2260 11880
rect 2500 11640 2590 11880
rect 2830 11640 2920 11880
rect 3160 11640 3250 11880
rect 3490 11640 3580 11880
rect 3820 11640 3910 11880
rect 4150 11640 4240 11880
rect 4480 11640 4570 11880
rect 4810 11640 4900 11880
rect 5140 11640 5230 11880
rect 5470 11640 5560 11880
rect 5800 11640 5890 11880
rect 6130 11640 6220 11880
rect 6460 11640 6550 11880
rect 6790 11640 6880 11880
rect 7120 11640 7290 11880
rect -5020 11550 7290 11640
rect -5020 11310 -4670 11550
rect -4430 11310 -4340 11550
rect -4100 11310 -4010 11550
rect -3770 11310 -3680 11550
rect -3440 11310 -3350 11550
rect -3110 11310 -3020 11550
rect -2780 11310 -2690 11550
rect -2450 11310 -2360 11550
rect -2120 11310 -2030 11550
rect -1790 11310 -1700 11550
rect -1460 11310 -1370 11550
rect -1130 11310 -1040 11550
rect -800 11310 -710 11550
rect -470 11310 -380 11550
rect -140 11310 -50 11550
rect 190 11310 280 11550
rect 520 11310 610 11550
rect 850 11310 940 11550
rect 1180 11310 1270 11550
rect 1510 11310 1600 11550
rect 1840 11310 1930 11550
rect 2170 11310 2260 11550
rect 2500 11310 2590 11550
rect 2830 11310 2920 11550
rect 3160 11310 3250 11550
rect 3490 11310 3580 11550
rect 3820 11310 3910 11550
rect 4150 11310 4240 11550
rect 4480 11310 4570 11550
rect 4810 11310 4900 11550
rect 5140 11310 5230 11550
rect 5470 11310 5560 11550
rect 5800 11310 5890 11550
rect 6130 11310 6220 11550
rect 6460 11310 6550 11550
rect 6790 11310 6880 11550
rect 7120 11310 7290 11550
rect -5020 11220 7290 11310
rect -5020 10980 -4670 11220
rect -4430 10980 -4340 11220
rect -4100 10980 -4010 11220
rect -3770 10980 -3680 11220
rect -3440 10980 -3350 11220
rect -3110 10980 -3020 11220
rect -2780 10980 -2690 11220
rect -2450 10980 -2360 11220
rect -2120 10980 -2030 11220
rect -1790 10980 -1700 11220
rect -1460 10980 -1370 11220
rect -1130 10980 -1040 11220
rect -800 10980 -710 11220
rect -470 10980 -380 11220
rect -140 10980 -50 11220
rect 190 10980 280 11220
rect 520 10980 610 11220
rect 850 10980 940 11220
rect 1180 10980 1270 11220
rect 1510 10980 1600 11220
rect 1840 10980 1930 11220
rect 2170 10980 2260 11220
rect 2500 10980 2590 11220
rect 2830 10980 2920 11220
rect 3160 10980 3250 11220
rect 3490 10980 3580 11220
rect 3820 10980 3910 11220
rect 4150 10980 4240 11220
rect 4480 10980 4570 11220
rect 4810 10980 4900 11220
rect 5140 10980 5230 11220
rect 5470 10980 5560 11220
rect 5800 10980 5890 11220
rect 6130 10980 6220 11220
rect 6460 10980 6550 11220
rect 6790 10980 6880 11220
rect 7120 10980 7290 11220
rect -5020 10890 7290 10980
rect -5020 10650 -4670 10890
rect -4430 10650 -4340 10890
rect -4100 10650 -4010 10890
rect -3770 10650 -3680 10890
rect -3440 10650 -3350 10890
rect -3110 10650 -3020 10890
rect -2780 10650 -2690 10890
rect -2450 10650 -2360 10890
rect -2120 10650 -2030 10890
rect -1790 10650 -1700 10890
rect -1460 10650 -1370 10890
rect -1130 10650 -1040 10890
rect -800 10650 -710 10890
rect -470 10650 -380 10890
rect -140 10650 -50 10890
rect 190 10650 280 10890
rect 520 10650 610 10890
rect 850 10650 940 10890
rect 1180 10650 1270 10890
rect 1510 10650 1600 10890
rect 1840 10650 1930 10890
rect 2170 10650 2260 10890
rect 2500 10650 2590 10890
rect 2830 10650 2920 10890
rect 3160 10650 3250 10890
rect 3490 10650 3580 10890
rect 3820 10650 3910 10890
rect 4150 10650 4240 10890
rect 4480 10650 4570 10890
rect 4810 10650 4900 10890
rect 5140 10650 5230 10890
rect 5470 10650 5560 10890
rect 5800 10650 5890 10890
rect 6130 10650 6220 10890
rect 6460 10650 6550 10890
rect 6790 10650 6880 10890
rect 7120 10650 7290 10890
rect -5020 10560 7290 10650
rect -5020 10320 -4670 10560
rect -4430 10320 -4340 10560
rect -4100 10320 -4010 10560
rect -3770 10320 -3680 10560
rect -3440 10320 -3350 10560
rect -3110 10320 -3020 10560
rect -2780 10320 -2690 10560
rect -2450 10320 -2360 10560
rect -2120 10320 -2030 10560
rect -1790 10320 -1700 10560
rect -1460 10320 -1370 10560
rect -1130 10320 -1040 10560
rect -800 10320 -710 10560
rect -470 10320 -380 10560
rect -140 10320 -50 10560
rect 190 10320 280 10560
rect 520 10320 610 10560
rect 850 10320 940 10560
rect 1180 10320 1270 10560
rect 1510 10320 1600 10560
rect 1840 10320 1930 10560
rect 2170 10320 2260 10560
rect 2500 10320 2590 10560
rect 2830 10320 2920 10560
rect 3160 10320 3250 10560
rect 3490 10320 3580 10560
rect 3820 10320 3910 10560
rect 4150 10320 4240 10560
rect 4480 10320 4570 10560
rect 4810 10320 4900 10560
rect 5140 10320 5230 10560
rect 5470 10320 5560 10560
rect 5800 10320 5890 10560
rect 6130 10320 6220 10560
rect 6460 10320 6550 10560
rect 6790 10320 6880 10560
rect 7120 10320 7290 10560
rect -5020 10230 7290 10320
rect -5020 9990 -4670 10230
rect -4430 9990 -4340 10230
rect -4100 9990 -4010 10230
rect -3770 9990 -3680 10230
rect -3440 9990 -3350 10230
rect -3110 9990 -3020 10230
rect -2780 9990 -2690 10230
rect -2450 9990 -2360 10230
rect -2120 9990 -2030 10230
rect -1790 9990 -1700 10230
rect -1460 9990 -1370 10230
rect -1130 9990 -1040 10230
rect -800 9990 -710 10230
rect -470 9990 -380 10230
rect -140 9990 -50 10230
rect 190 9990 280 10230
rect 520 9990 610 10230
rect 850 9990 940 10230
rect 1180 9990 1270 10230
rect 1510 9990 1600 10230
rect 1840 9990 1930 10230
rect 2170 9990 2260 10230
rect 2500 9990 2590 10230
rect 2830 9990 2920 10230
rect 3160 9990 3250 10230
rect 3490 9990 3580 10230
rect 3820 9990 3910 10230
rect 4150 9990 4240 10230
rect 4480 9990 4570 10230
rect 4810 9990 4900 10230
rect 5140 9990 5230 10230
rect 5470 9990 5560 10230
rect 5800 9990 5890 10230
rect 6130 9990 6220 10230
rect 6460 9990 6550 10230
rect 6790 9990 6880 10230
rect 7120 9990 7290 10230
rect -5020 9900 7290 9990
rect -5020 9660 -4670 9900
rect -4430 9660 -4340 9900
rect -4100 9660 -4010 9900
rect -3770 9660 -3680 9900
rect -3440 9660 -3350 9900
rect -3110 9660 -3020 9900
rect -2780 9660 -2690 9900
rect -2450 9660 -2360 9900
rect -2120 9660 -2030 9900
rect -1790 9660 -1700 9900
rect -1460 9660 -1370 9900
rect -1130 9660 -1040 9900
rect -800 9660 -710 9900
rect -470 9660 -380 9900
rect -140 9660 -50 9900
rect 190 9660 280 9900
rect 520 9660 610 9900
rect 850 9660 940 9900
rect 1180 9660 1270 9900
rect 1510 9660 1600 9900
rect 1840 9660 1930 9900
rect 2170 9660 2260 9900
rect 2500 9660 2590 9900
rect 2830 9660 2920 9900
rect 3160 9660 3250 9900
rect 3490 9660 3580 9900
rect 3820 9660 3910 9900
rect 4150 9660 4240 9900
rect 4480 9660 4570 9900
rect 4810 9660 4900 9900
rect 5140 9660 5230 9900
rect 5470 9660 5560 9900
rect 5800 9660 5890 9900
rect 6130 9660 6220 9900
rect 6460 9660 6550 9900
rect 6790 9660 6880 9900
rect 7120 9660 7290 9900
rect -5020 9570 7290 9660
rect -5020 9330 -4670 9570
rect -4430 9330 -4340 9570
rect -4100 9330 -4010 9570
rect -3770 9330 -3680 9570
rect -3440 9330 -3350 9570
rect -3110 9330 -3020 9570
rect -2780 9330 -2690 9570
rect -2450 9330 -2360 9570
rect -2120 9330 -2030 9570
rect -1790 9330 -1700 9570
rect -1460 9330 -1370 9570
rect -1130 9330 -1040 9570
rect -800 9330 -710 9570
rect -470 9330 -380 9570
rect -140 9330 -50 9570
rect 190 9330 280 9570
rect 520 9330 610 9570
rect 850 9330 940 9570
rect 1180 9330 1270 9570
rect 1510 9330 1600 9570
rect 1840 9330 1930 9570
rect 2170 9330 2260 9570
rect 2500 9330 2590 9570
rect 2830 9330 2920 9570
rect 3160 9330 3250 9570
rect 3490 9330 3580 9570
rect 3820 9330 3910 9570
rect 4150 9330 4240 9570
rect 4480 9330 4570 9570
rect 4810 9330 4900 9570
rect 5140 9330 5230 9570
rect 5470 9330 5560 9570
rect 5800 9330 5890 9570
rect 6130 9330 6220 9570
rect 6460 9330 6550 9570
rect 6790 9330 6880 9570
rect 7120 9330 7290 9570
rect -5020 9240 7290 9330
rect -5020 9000 -4670 9240
rect -4430 9000 -4340 9240
rect -4100 9000 -4010 9240
rect -3770 9000 -3680 9240
rect -3440 9000 -3350 9240
rect -3110 9000 -3020 9240
rect -2780 9000 -2690 9240
rect -2450 9000 -2360 9240
rect -2120 9000 -2030 9240
rect -1790 9000 -1700 9240
rect -1460 9000 -1370 9240
rect -1130 9000 -1040 9240
rect -800 9000 -710 9240
rect -470 9000 -380 9240
rect -140 9000 -50 9240
rect 190 9000 280 9240
rect 520 9000 610 9240
rect 850 9000 940 9240
rect 1180 9000 1270 9240
rect 1510 9000 1600 9240
rect 1840 9000 1930 9240
rect 2170 9000 2260 9240
rect 2500 9000 2590 9240
rect 2830 9000 2920 9240
rect 3160 9000 3250 9240
rect 3490 9000 3580 9240
rect 3820 9000 3910 9240
rect 4150 9000 4240 9240
rect 4480 9000 4570 9240
rect 4810 9000 4900 9240
rect 5140 9000 5230 9240
rect 5470 9000 5560 9240
rect 5800 9000 5890 9240
rect 6130 9000 6220 9240
rect 6460 9000 6550 9240
rect 6790 9000 6880 9240
rect 7120 9000 7290 9240
rect -5020 8830 7290 9000
rect 7610 21140 7880 21300
rect 7610 20790 19920 21140
rect 7610 20550 7780 20790
rect 8020 20550 8110 20790
rect 8350 20550 8440 20790
rect 8680 20550 8770 20790
rect 9010 20550 9100 20790
rect 9340 20550 9430 20790
rect 9670 20550 9760 20790
rect 10000 20550 10090 20790
rect 10330 20550 10420 20790
rect 10660 20550 10750 20790
rect 10990 20550 11080 20790
rect 11320 20550 11410 20790
rect 11650 20550 11740 20790
rect 11980 20550 12070 20790
rect 12310 20550 12400 20790
rect 12640 20550 12730 20790
rect 12970 20550 13060 20790
rect 13300 20550 13390 20790
rect 13630 20550 13720 20790
rect 13960 20550 14050 20790
rect 14290 20550 14380 20790
rect 14620 20550 14710 20790
rect 14950 20550 15040 20790
rect 15280 20550 15370 20790
rect 15610 20550 15700 20790
rect 15940 20550 16030 20790
rect 16270 20550 16360 20790
rect 16600 20550 16690 20790
rect 16930 20550 17020 20790
rect 17260 20550 17350 20790
rect 17590 20550 17680 20790
rect 17920 20550 18010 20790
rect 18250 20550 18340 20790
rect 18580 20550 18670 20790
rect 18910 20550 19000 20790
rect 19240 20550 19330 20790
rect 19570 20550 19920 20790
rect 7610 20460 19920 20550
rect 7610 20220 7780 20460
rect 8020 20220 8110 20460
rect 8350 20220 8440 20460
rect 8680 20220 8770 20460
rect 9010 20220 9100 20460
rect 9340 20220 9430 20460
rect 9670 20220 9760 20460
rect 10000 20220 10090 20460
rect 10330 20220 10420 20460
rect 10660 20220 10750 20460
rect 10990 20220 11080 20460
rect 11320 20220 11410 20460
rect 11650 20220 11740 20460
rect 11980 20220 12070 20460
rect 12310 20220 12400 20460
rect 12640 20220 12730 20460
rect 12970 20220 13060 20460
rect 13300 20220 13390 20460
rect 13630 20220 13720 20460
rect 13960 20220 14050 20460
rect 14290 20220 14380 20460
rect 14620 20220 14710 20460
rect 14950 20220 15040 20460
rect 15280 20220 15370 20460
rect 15610 20220 15700 20460
rect 15940 20220 16030 20460
rect 16270 20220 16360 20460
rect 16600 20220 16690 20460
rect 16930 20220 17020 20460
rect 17260 20220 17350 20460
rect 17590 20220 17680 20460
rect 17920 20220 18010 20460
rect 18250 20220 18340 20460
rect 18580 20220 18670 20460
rect 18910 20220 19000 20460
rect 19240 20220 19330 20460
rect 19570 20220 19920 20460
rect 7610 20130 19920 20220
rect 7610 19890 7780 20130
rect 8020 19890 8110 20130
rect 8350 19890 8440 20130
rect 8680 19890 8770 20130
rect 9010 19890 9100 20130
rect 9340 19890 9430 20130
rect 9670 19890 9760 20130
rect 10000 19890 10090 20130
rect 10330 19890 10420 20130
rect 10660 19890 10750 20130
rect 10990 19890 11080 20130
rect 11320 19890 11410 20130
rect 11650 19890 11740 20130
rect 11980 19890 12070 20130
rect 12310 19890 12400 20130
rect 12640 19890 12730 20130
rect 12970 19890 13060 20130
rect 13300 19890 13390 20130
rect 13630 19890 13720 20130
rect 13960 19890 14050 20130
rect 14290 19890 14380 20130
rect 14620 19890 14710 20130
rect 14950 19890 15040 20130
rect 15280 19890 15370 20130
rect 15610 19890 15700 20130
rect 15940 19890 16030 20130
rect 16270 19890 16360 20130
rect 16600 19890 16690 20130
rect 16930 19890 17020 20130
rect 17260 19890 17350 20130
rect 17590 19890 17680 20130
rect 17920 19890 18010 20130
rect 18250 19890 18340 20130
rect 18580 19890 18670 20130
rect 18910 19890 19000 20130
rect 19240 19890 19330 20130
rect 19570 19890 19920 20130
rect 7610 19800 19920 19890
rect 7610 19560 7780 19800
rect 8020 19560 8110 19800
rect 8350 19560 8440 19800
rect 8680 19560 8770 19800
rect 9010 19560 9100 19800
rect 9340 19560 9430 19800
rect 9670 19560 9760 19800
rect 10000 19560 10090 19800
rect 10330 19560 10420 19800
rect 10660 19560 10750 19800
rect 10990 19560 11080 19800
rect 11320 19560 11410 19800
rect 11650 19560 11740 19800
rect 11980 19560 12070 19800
rect 12310 19560 12400 19800
rect 12640 19560 12730 19800
rect 12970 19560 13060 19800
rect 13300 19560 13390 19800
rect 13630 19560 13720 19800
rect 13960 19560 14050 19800
rect 14290 19560 14380 19800
rect 14620 19560 14710 19800
rect 14950 19560 15040 19800
rect 15280 19560 15370 19800
rect 15610 19560 15700 19800
rect 15940 19560 16030 19800
rect 16270 19560 16360 19800
rect 16600 19560 16690 19800
rect 16930 19560 17020 19800
rect 17260 19560 17350 19800
rect 17590 19560 17680 19800
rect 17920 19560 18010 19800
rect 18250 19560 18340 19800
rect 18580 19560 18670 19800
rect 18910 19560 19000 19800
rect 19240 19560 19330 19800
rect 19570 19560 19920 19800
rect 7610 19470 19920 19560
rect 7610 19230 7780 19470
rect 8020 19230 8110 19470
rect 8350 19230 8440 19470
rect 8680 19230 8770 19470
rect 9010 19230 9100 19470
rect 9340 19230 9430 19470
rect 9670 19230 9760 19470
rect 10000 19230 10090 19470
rect 10330 19230 10420 19470
rect 10660 19230 10750 19470
rect 10990 19230 11080 19470
rect 11320 19230 11410 19470
rect 11650 19230 11740 19470
rect 11980 19230 12070 19470
rect 12310 19230 12400 19470
rect 12640 19230 12730 19470
rect 12970 19230 13060 19470
rect 13300 19230 13390 19470
rect 13630 19230 13720 19470
rect 13960 19230 14050 19470
rect 14290 19230 14380 19470
rect 14620 19230 14710 19470
rect 14950 19230 15040 19470
rect 15280 19230 15370 19470
rect 15610 19230 15700 19470
rect 15940 19230 16030 19470
rect 16270 19230 16360 19470
rect 16600 19230 16690 19470
rect 16930 19230 17020 19470
rect 17260 19230 17350 19470
rect 17590 19230 17680 19470
rect 17920 19230 18010 19470
rect 18250 19230 18340 19470
rect 18580 19230 18670 19470
rect 18910 19230 19000 19470
rect 19240 19230 19330 19470
rect 19570 19230 19920 19470
rect 7610 19140 19920 19230
rect 7610 18900 7780 19140
rect 8020 18900 8110 19140
rect 8350 18900 8440 19140
rect 8680 18900 8770 19140
rect 9010 18900 9100 19140
rect 9340 18900 9430 19140
rect 9670 18900 9760 19140
rect 10000 18900 10090 19140
rect 10330 18900 10420 19140
rect 10660 18900 10750 19140
rect 10990 18900 11080 19140
rect 11320 18900 11410 19140
rect 11650 18900 11740 19140
rect 11980 18900 12070 19140
rect 12310 18900 12400 19140
rect 12640 18900 12730 19140
rect 12970 18900 13060 19140
rect 13300 18900 13390 19140
rect 13630 18900 13720 19140
rect 13960 18900 14050 19140
rect 14290 18900 14380 19140
rect 14620 18900 14710 19140
rect 14950 18900 15040 19140
rect 15280 18900 15370 19140
rect 15610 18900 15700 19140
rect 15940 18900 16030 19140
rect 16270 18900 16360 19140
rect 16600 18900 16690 19140
rect 16930 18900 17020 19140
rect 17260 18900 17350 19140
rect 17590 18900 17680 19140
rect 17920 18900 18010 19140
rect 18250 18900 18340 19140
rect 18580 18900 18670 19140
rect 18910 18900 19000 19140
rect 19240 18900 19330 19140
rect 19570 18900 19920 19140
rect 7610 18810 19920 18900
rect 7610 18570 7780 18810
rect 8020 18570 8110 18810
rect 8350 18570 8440 18810
rect 8680 18570 8770 18810
rect 9010 18570 9100 18810
rect 9340 18570 9430 18810
rect 9670 18570 9760 18810
rect 10000 18570 10090 18810
rect 10330 18570 10420 18810
rect 10660 18570 10750 18810
rect 10990 18570 11080 18810
rect 11320 18570 11410 18810
rect 11650 18570 11740 18810
rect 11980 18570 12070 18810
rect 12310 18570 12400 18810
rect 12640 18570 12730 18810
rect 12970 18570 13060 18810
rect 13300 18570 13390 18810
rect 13630 18570 13720 18810
rect 13960 18570 14050 18810
rect 14290 18570 14380 18810
rect 14620 18570 14710 18810
rect 14950 18570 15040 18810
rect 15280 18570 15370 18810
rect 15610 18570 15700 18810
rect 15940 18570 16030 18810
rect 16270 18570 16360 18810
rect 16600 18570 16690 18810
rect 16930 18570 17020 18810
rect 17260 18570 17350 18810
rect 17590 18570 17680 18810
rect 17920 18570 18010 18810
rect 18250 18570 18340 18810
rect 18580 18570 18670 18810
rect 18910 18570 19000 18810
rect 19240 18570 19330 18810
rect 19570 18570 19920 18810
rect 7610 18480 19920 18570
rect 7610 18240 7780 18480
rect 8020 18240 8110 18480
rect 8350 18240 8440 18480
rect 8680 18240 8770 18480
rect 9010 18240 9100 18480
rect 9340 18240 9430 18480
rect 9670 18240 9760 18480
rect 10000 18240 10090 18480
rect 10330 18240 10420 18480
rect 10660 18240 10750 18480
rect 10990 18240 11080 18480
rect 11320 18240 11410 18480
rect 11650 18240 11740 18480
rect 11980 18240 12070 18480
rect 12310 18240 12400 18480
rect 12640 18240 12730 18480
rect 12970 18240 13060 18480
rect 13300 18240 13390 18480
rect 13630 18240 13720 18480
rect 13960 18240 14050 18480
rect 14290 18240 14380 18480
rect 14620 18240 14710 18480
rect 14950 18240 15040 18480
rect 15280 18240 15370 18480
rect 15610 18240 15700 18480
rect 15940 18240 16030 18480
rect 16270 18240 16360 18480
rect 16600 18240 16690 18480
rect 16930 18240 17020 18480
rect 17260 18240 17350 18480
rect 17590 18240 17680 18480
rect 17920 18240 18010 18480
rect 18250 18240 18340 18480
rect 18580 18240 18670 18480
rect 18910 18240 19000 18480
rect 19240 18240 19330 18480
rect 19570 18240 19920 18480
rect 7610 18150 19920 18240
rect 7610 17910 7780 18150
rect 8020 17910 8110 18150
rect 8350 17910 8440 18150
rect 8680 17910 8770 18150
rect 9010 17910 9100 18150
rect 9340 17910 9430 18150
rect 9670 17910 9760 18150
rect 10000 17910 10090 18150
rect 10330 17910 10420 18150
rect 10660 17910 10750 18150
rect 10990 17910 11080 18150
rect 11320 17910 11410 18150
rect 11650 17910 11740 18150
rect 11980 17910 12070 18150
rect 12310 17910 12400 18150
rect 12640 17910 12730 18150
rect 12970 17910 13060 18150
rect 13300 17910 13390 18150
rect 13630 17910 13720 18150
rect 13960 17910 14050 18150
rect 14290 17910 14380 18150
rect 14620 17910 14710 18150
rect 14950 17910 15040 18150
rect 15280 17910 15370 18150
rect 15610 17910 15700 18150
rect 15940 17910 16030 18150
rect 16270 17910 16360 18150
rect 16600 17910 16690 18150
rect 16930 17910 17020 18150
rect 17260 17910 17350 18150
rect 17590 17910 17680 18150
rect 17920 17910 18010 18150
rect 18250 17910 18340 18150
rect 18580 17910 18670 18150
rect 18910 17910 19000 18150
rect 19240 17910 19330 18150
rect 19570 17910 19920 18150
rect 7610 17820 19920 17910
rect 7610 17580 7780 17820
rect 8020 17580 8110 17820
rect 8350 17580 8440 17820
rect 8680 17580 8770 17820
rect 9010 17580 9100 17820
rect 9340 17580 9430 17820
rect 9670 17580 9760 17820
rect 10000 17580 10090 17820
rect 10330 17580 10420 17820
rect 10660 17580 10750 17820
rect 10990 17580 11080 17820
rect 11320 17580 11410 17820
rect 11650 17580 11740 17820
rect 11980 17580 12070 17820
rect 12310 17580 12400 17820
rect 12640 17580 12730 17820
rect 12970 17580 13060 17820
rect 13300 17580 13390 17820
rect 13630 17580 13720 17820
rect 13960 17580 14050 17820
rect 14290 17580 14380 17820
rect 14620 17580 14710 17820
rect 14950 17580 15040 17820
rect 15280 17580 15370 17820
rect 15610 17580 15700 17820
rect 15940 17580 16030 17820
rect 16270 17580 16360 17820
rect 16600 17580 16690 17820
rect 16930 17580 17020 17820
rect 17260 17580 17350 17820
rect 17590 17580 17680 17820
rect 17920 17580 18010 17820
rect 18250 17580 18340 17820
rect 18580 17580 18670 17820
rect 18910 17580 19000 17820
rect 19240 17580 19330 17820
rect 19570 17580 19920 17820
rect 7610 17490 19920 17580
rect 7610 17250 7780 17490
rect 8020 17250 8110 17490
rect 8350 17250 8440 17490
rect 8680 17250 8770 17490
rect 9010 17250 9100 17490
rect 9340 17250 9430 17490
rect 9670 17250 9760 17490
rect 10000 17250 10090 17490
rect 10330 17250 10420 17490
rect 10660 17250 10750 17490
rect 10990 17250 11080 17490
rect 11320 17250 11410 17490
rect 11650 17250 11740 17490
rect 11980 17250 12070 17490
rect 12310 17250 12400 17490
rect 12640 17250 12730 17490
rect 12970 17250 13060 17490
rect 13300 17250 13390 17490
rect 13630 17250 13720 17490
rect 13960 17250 14050 17490
rect 14290 17250 14380 17490
rect 14620 17250 14710 17490
rect 14950 17250 15040 17490
rect 15280 17250 15370 17490
rect 15610 17250 15700 17490
rect 15940 17250 16030 17490
rect 16270 17250 16360 17490
rect 16600 17250 16690 17490
rect 16930 17250 17020 17490
rect 17260 17250 17350 17490
rect 17590 17250 17680 17490
rect 17920 17250 18010 17490
rect 18250 17250 18340 17490
rect 18580 17250 18670 17490
rect 18910 17250 19000 17490
rect 19240 17250 19330 17490
rect 19570 17250 19920 17490
rect 7610 17160 19920 17250
rect 7610 16920 7780 17160
rect 8020 16920 8110 17160
rect 8350 16920 8440 17160
rect 8680 16920 8770 17160
rect 9010 16920 9100 17160
rect 9340 16920 9430 17160
rect 9670 16920 9760 17160
rect 10000 16920 10090 17160
rect 10330 16920 10420 17160
rect 10660 16920 10750 17160
rect 10990 16920 11080 17160
rect 11320 16920 11410 17160
rect 11650 16920 11740 17160
rect 11980 16920 12070 17160
rect 12310 16920 12400 17160
rect 12640 16920 12730 17160
rect 12970 16920 13060 17160
rect 13300 16920 13390 17160
rect 13630 16920 13720 17160
rect 13960 16920 14050 17160
rect 14290 16920 14380 17160
rect 14620 16920 14710 17160
rect 14950 16920 15040 17160
rect 15280 16920 15370 17160
rect 15610 16920 15700 17160
rect 15940 16920 16030 17160
rect 16270 16920 16360 17160
rect 16600 16920 16690 17160
rect 16930 16920 17020 17160
rect 17260 16920 17350 17160
rect 17590 16920 17680 17160
rect 17920 16920 18010 17160
rect 18250 16920 18340 17160
rect 18580 16920 18670 17160
rect 18910 16920 19000 17160
rect 19240 16920 19330 17160
rect 19570 16920 19920 17160
rect 7610 16830 19920 16920
rect 7610 16590 7780 16830
rect 8020 16590 8110 16830
rect 8350 16590 8440 16830
rect 8680 16590 8770 16830
rect 9010 16590 9100 16830
rect 9340 16590 9430 16830
rect 9670 16590 9760 16830
rect 10000 16590 10090 16830
rect 10330 16590 10420 16830
rect 10660 16590 10750 16830
rect 10990 16590 11080 16830
rect 11320 16590 11410 16830
rect 11650 16590 11740 16830
rect 11980 16590 12070 16830
rect 12310 16590 12400 16830
rect 12640 16590 12730 16830
rect 12970 16590 13060 16830
rect 13300 16590 13390 16830
rect 13630 16590 13720 16830
rect 13960 16590 14050 16830
rect 14290 16590 14380 16830
rect 14620 16590 14710 16830
rect 14950 16590 15040 16830
rect 15280 16590 15370 16830
rect 15610 16590 15700 16830
rect 15940 16590 16030 16830
rect 16270 16590 16360 16830
rect 16600 16590 16690 16830
rect 16930 16590 17020 16830
rect 17260 16590 17350 16830
rect 17590 16590 17680 16830
rect 17920 16590 18010 16830
rect 18250 16590 18340 16830
rect 18580 16590 18670 16830
rect 18910 16590 19000 16830
rect 19240 16590 19330 16830
rect 19570 16590 19920 16830
rect 7610 16500 19920 16590
rect 7610 16260 7780 16500
rect 8020 16260 8110 16500
rect 8350 16260 8440 16500
rect 8680 16260 8770 16500
rect 9010 16260 9100 16500
rect 9340 16260 9430 16500
rect 9670 16260 9760 16500
rect 10000 16260 10090 16500
rect 10330 16260 10420 16500
rect 10660 16260 10750 16500
rect 10990 16260 11080 16500
rect 11320 16260 11410 16500
rect 11650 16260 11740 16500
rect 11980 16260 12070 16500
rect 12310 16260 12400 16500
rect 12640 16260 12730 16500
rect 12970 16260 13060 16500
rect 13300 16260 13390 16500
rect 13630 16260 13720 16500
rect 13960 16260 14050 16500
rect 14290 16260 14380 16500
rect 14620 16260 14710 16500
rect 14950 16260 15040 16500
rect 15280 16260 15370 16500
rect 15610 16260 15700 16500
rect 15940 16260 16030 16500
rect 16270 16260 16360 16500
rect 16600 16260 16690 16500
rect 16930 16260 17020 16500
rect 17260 16260 17350 16500
rect 17590 16260 17680 16500
rect 17920 16260 18010 16500
rect 18250 16260 18340 16500
rect 18580 16260 18670 16500
rect 18910 16260 19000 16500
rect 19240 16260 19330 16500
rect 19570 16260 19920 16500
rect 7610 16170 19920 16260
rect 7610 15930 7780 16170
rect 8020 15930 8110 16170
rect 8350 15930 8440 16170
rect 8680 15930 8770 16170
rect 9010 15930 9100 16170
rect 9340 15930 9430 16170
rect 9670 15930 9760 16170
rect 10000 15930 10090 16170
rect 10330 15930 10420 16170
rect 10660 15930 10750 16170
rect 10990 15930 11080 16170
rect 11320 15930 11410 16170
rect 11650 15930 11740 16170
rect 11980 15930 12070 16170
rect 12310 15930 12400 16170
rect 12640 15930 12730 16170
rect 12970 15930 13060 16170
rect 13300 15930 13390 16170
rect 13630 15930 13720 16170
rect 13960 15930 14050 16170
rect 14290 15930 14380 16170
rect 14620 15930 14710 16170
rect 14950 15930 15040 16170
rect 15280 15930 15370 16170
rect 15610 15930 15700 16170
rect 15940 15930 16030 16170
rect 16270 15930 16360 16170
rect 16600 15930 16690 16170
rect 16930 15930 17020 16170
rect 17260 15930 17350 16170
rect 17590 15930 17680 16170
rect 17920 15930 18010 16170
rect 18250 15930 18340 16170
rect 18580 15930 18670 16170
rect 18910 15930 19000 16170
rect 19240 15930 19330 16170
rect 19570 15930 19920 16170
rect 7610 15840 19920 15930
rect 7610 15600 7780 15840
rect 8020 15600 8110 15840
rect 8350 15600 8440 15840
rect 8680 15600 8770 15840
rect 9010 15600 9100 15840
rect 9340 15600 9430 15840
rect 9670 15600 9760 15840
rect 10000 15600 10090 15840
rect 10330 15600 10420 15840
rect 10660 15600 10750 15840
rect 10990 15600 11080 15840
rect 11320 15600 11410 15840
rect 11650 15600 11740 15840
rect 11980 15600 12070 15840
rect 12310 15600 12400 15840
rect 12640 15600 12730 15840
rect 12970 15600 13060 15840
rect 13300 15600 13390 15840
rect 13630 15600 13720 15840
rect 13960 15600 14050 15840
rect 14290 15600 14380 15840
rect 14620 15600 14710 15840
rect 14950 15600 15040 15840
rect 15280 15600 15370 15840
rect 15610 15600 15700 15840
rect 15940 15600 16030 15840
rect 16270 15600 16360 15840
rect 16600 15600 16690 15840
rect 16930 15600 17020 15840
rect 17260 15600 17350 15840
rect 17590 15600 17680 15840
rect 17920 15600 18010 15840
rect 18250 15600 18340 15840
rect 18580 15600 18670 15840
rect 18910 15600 19000 15840
rect 19240 15600 19330 15840
rect 19570 15600 19920 15840
rect 7610 15510 19920 15600
rect 7610 15270 7780 15510
rect 8020 15270 8110 15510
rect 8350 15270 8440 15510
rect 8680 15270 8770 15510
rect 9010 15270 9100 15510
rect 9340 15270 9430 15510
rect 9670 15270 9760 15510
rect 10000 15270 10090 15510
rect 10330 15270 10420 15510
rect 10660 15270 10750 15510
rect 10990 15270 11080 15510
rect 11320 15270 11410 15510
rect 11650 15270 11740 15510
rect 11980 15270 12070 15510
rect 12310 15270 12400 15510
rect 12640 15270 12730 15510
rect 12970 15270 13060 15510
rect 13300 15270 13390 15510
rect 13630 15270 13720 15510
rect 13960 15270 14050 15510
rect 14290 15270 14380 15510
rect 14620 15270 14710 15510
rect 14950 15270 15040 15510
rect 15280 15270 15370 15510
rect 15610 15270 15700 15510
rect 15940 15270 16030 15510
rect 16270 15270 16360 15510
rect 16600 15270 16690 15510
rect 16930 15270 17020 15510
rect 17260 15270 17350 15510
rect 17590 15270 17680 15510
rect 17920 15270 18010 15510
rect 18250 15270 18340 15510
rect 18580 15270 18670 15510
rect 18910 15270 19000 15510
rect 19240 15270 19330 15510
rect 19570 15270 19920 15510
rect 7610 15180 19920 15270
rect 7610 14940 7780 15180
rect 8020 14940 8110 15180
rect 8350 14940 8440 15180
rect 8680 14940 8770 15180
rect 9010 14940 9100 15180
rect 9340 14940 9430 15180
rect 9670 14940 9760 15180
rect 10000 14940 10090 15180
rect 10330 14940 10420 15180
rect 10660 14940 10750 15180
rect 10990 14940 11080 15180
rect 11320 14940 11410 15180
rect 11650 14940 11740 15180
rect 11980 14940 12070 15180
rect 12310 14940 12400 15180
rect 12640 14940 12730 15180
rect 12970 14940 13060 15180
rect 13300 14940 13390 15180
rect 13630 14940 13720 15180
rect 13960 14940 14050 15180
rect 14290 14940 14380 15180
rect 14620 14940 14710 15180
rect 14950 14940 15040 15180
rect 15280 14940 15370 15180
rect 15610 14940 15700 15180
rect 15940 14940 16030 15180
rect 16270 14940 16360 15180
rect 16600 14940 16690 15180
rect 16930 14940 17020 15180
rect 17260 14940 17350 15180
rect 17590 14940 17680 15180
rect 17920 14940 18010 15180
rect 18250 14940 18340 15180
rect 18580 14940 18670 15180
rect 18910 14940 19000 15180
rect 19240 14940 19330 15180
rect 19570 14940 19920 15180
rect 7610 14850 19920 14940
rect 7610 14610 7780 14850
rect 8020 14610 8110 14850
rect 8350 14610 8440 14850
rect 8680 14610 8770 14850
rect 9010 14610 9100 14850
rect 9340 14610 9430 14850
rect 9670 14610 9760 14850
rect 10000 14610 10090 14850
rect 10330 14610 10420 14850
rect 10660 14610 10750 14850
rect 10990 14610 11080 14850
rect 11320 14610 11410 14850
rect 11650 14610 11740 14850
rect 11980 14610 12070 14850
rect 12310 14610 12400 14850
rect 12640 14610 12730 14850
rect 12970 14610 13060 14850
rect 13300 14610 13390 14850
rect 13630 14610 13720 14850
rect 13960 14610 14050 14850
rect 14290 14610 14380 14850
rect 14620 14610 14710 14850
rect 14950 14610 15040 14850
rect 15280 14610 15370 14850
rect 15610 14610 15700 14850
rect 15940 14610 16030 14850
rect 16270 14610 16360 14850
rect 16600 14610 16690 14850
rect 16930 14610 17020 14850
rect 17260 14610 17350 14850
rect 17590 14610 17680 14850
rect 17920 14610 18010 14850
rect 18250 14610 18340 14850
rect 18580 14610 18670 14850
rect 18910 14610 19000 14850
rect 19240 14610 19330 14850
rect 19570 14610 19920 14850
rect 7610 14520 19920 14610
rect 7610 14280 7780 14520
rect 8020 14280 8110 14520
rect 8350 14280 8440 14520
rect 8680 14280 8770 14520
rect 9010 14280 9100 14520
rect 9340 14280 9430 14520
rect 9670 14280 9760 14520
rect 10000 14280 10090 14520
rect 10330 14280 10420 14520
rect 10660 14280 10750 14520
rect 10990 14280 11080 14520
rect 11320 14280 11410 14520
rect 11650 14280 11740 14520
rect 11980 14280 12070 14520
rect 12310 14280 12400 14520
rect 12640 14280 12730 14520
rect 12970 14280 13060 14520
rect 13300 14280 13390 14520
rect 13630 14280 13720 14520
rect 13960 14280 14050 14520
rect 14290 14280 14380 14520
rect 14620 14280 14710 14520
rect 14950 14280 15040 14520
rect 15280 14280 15370 14520
rect 15610 14280 15700 14520
rect 15940 14280 16030 14520
rect 16270 14280 16360 14520
rect 16600 14280 16690 14520
rect 16930 14280 17020 14520
rect 17260 14280 17350 14520
rect 17590 14280 17680 14520
rect 17920 14280 18010 14520
rect 18250 14280 18340 14520
rect 18580 14280 18670 14520
rect 18910 14280 19000 14520
rect 19240 14280 19330 14520
rect 19570 14280 19920 14520
rect 7610 14190 19920 14280
rect 7610 13950 7780 14190
rect 8020 13950 8110 14190
rect 8350 13950 8440 14190
rect 8680 13950 8770 14190
rect 9010 13950 9100 14190
rect 9340 13950 9430 14190
rect 9670 13950 9760 14190
rect 10000 13950 10090 14190
rect 10330 13950 10420 14190
rect 10660 13950 10750 14190
rect 10990 13950 11080 14190
rect 11320 13950 11410 14190
rect 11650 13950 11740 14190
rect 11980 13950 12070 14190
rect 12310 13950 12400 14190
rect 12640 13950 12730 14190
rect 12970 13950 13060 14190
rect 13300 13950 13390 14190
rect 13630 13950 13720 14190
rect 13960 13950 14050 14190
rect 14290 13950 14380 14190
rect 14620 13950 14710 14190
rect 14950 13950 15040 14190
rect 15280 13950 15370 14190
rect 15610 13950 15700 14190
rect 15940 13950 16030 14190
rect 16270 13950 16360 14190
rect 16600 13950 16690 14190
rect 16930 13950 17020 14190
rect 17260 13950 17350 14190
rect 17590 13950 17680 14190
rect 17920 13950 18010 14190
rect 18250 13950 18340 14190
rect 18580 13950 18670 14190
rect 18910 13950 19000 14190
rect 19240 13950 19330 14190
rect 19570 13950 19920 14190
rect 7610 13860 19920 13950
rect 7610 13620 7780 13860
rect 8020 13620 8110 13860
rect 8350 13620 8440 13860
rect 8680 13620 8770 13860
rect 9010 13620 9100 13860
rect 9340 13620 9430 13860
rect 9670 13620 9760 13860
rect 10000 13620 10090 13860
rect 10330 13620 10420 13860
rect 10660 13620 10750 13860
rect 10990 13620 11080 13860
rect 11320 13620 11410 13860
rect 11650 13620 11740 13860
rect 11980 13620 12070 13860
rect 12310 13620 12400 13860
rect 12640 13620 12730 13860
rect 12970 13620 13060 13860
rect 13300 13620 13390 13860
rect 13630 13620 13720 13860
rect 13960 13620 14050 13860
rect 14290 13620 14380 13860
rect 14620 13620 14710 13860
rect 14950 13620 15040 13860
rect 15280 13620 15370 13860
rect 15610 13620 15700 13860
rect 15940 13620 16030 13860
rect 16270 13620 16360 13860
rect 16600 13620 16690 13860
rect 16930 13620 17020 13860
rect 17260 13620 17350 13860
rect 17590 13620 17680 13860
rect 17920 13620 18010 13860
rect 18250 13620 18340 13860
rect 18580 13620 18670 13860
rect 18910 13620 19000 13860
rect 19240 13620 19330 13860
rect 19570 13620 19920 13860
rect 7610 13530 19920 13620
rect 7610 13290 7780 13530
rect 8020 13290 8110 13530
rect 8350 13290 8440 13530
rect 8680 13290 8770 13530
rect 9010 13290 9100 13530
rect 9340 13290 9430 13530
rect 9670 13290 9760 13530
rect 10000 13290 10090 13530
rect 10330 13290 10420 13530
rect 10660 13290 10750 13530
rect 10990 13290 11080 13530
rect 11320 13290 11410 13530
rect 11650 13290 11740 13530
rect 11980 13290 12070 13530
rect 12310 13290 12400 13530
rect 12640 13290 12730 13530
rect 12970 13290 13060 13530
rect 13300 13290 13390 13530
rect 13630 13290 13720 13530
rect 13960 13290 14050 13530
rect 14290 13290 14380 13530
rect 14620 13290 14710 13530
rect 14950 13290 15040 13530
rect 15280 13290 15370 13530
rect 15610 13290 15700 13530
rect 15940 13290 16030 13530
rect 16270 13290 16360 13530
rect 16600 13290 16690 13530
rect 16930 13290 17020 13530
rect 17260 13290 17350 13530
rect 17590 13290 17680 13530
rect 17920 13290 18010 13530
rect 18250 13290 18340 13530
rect 18580 13290 18670 13530
rect 18910 13290 19000 13530
rect 19240 13290 19330 13530
rect 19570 13290 19920 13530
rect 7610 13200 19920 13290
rect 7610 12960 7780 13200
rect 8020 12960 8110 13200
rect 8350 12960 8440 13200
rect 8680 12960 8770 13200
rect 9010 12960 9100 13200
rect 9340 12960 9430 13200
rect 9670 12960 9760 13200
rect 10000 12960 10090 13200
rect 10330 12960 10420 13200
rect 10660 12960 10750 13200
rect 10990 12960 11080 13200
rect 11320 12960 11410 13200
rect 11650 12960 11740 13200
rect 11980 12960 12070 13200
rect 12310 12960 12400 13200
rect 12640 12960 12730 13200
rect 12970 12960 13060 13200
rect 13300 12960 13390 13200
rect 13630 12960 13720 13200
rect 13960 12960 14050 13200
rect 14290 12960 14380 13200
rect 14620 12960 14710 13200
rect 14950 12960 15040 13200
rect 15280 12960 15370 13200
rect 15610 12960 15700 13200
rect 15940 12960 16030 13200
rect 16270 12960 16360 13200
rect 16600 12960 16690 13200
rect 16930 12960 17020 13200
rect 17260 12960 17350 13200
rect 17590 12960 17680 13200
rect 17920 12960 18010 13200
rect 18250 12960 18340 13200
rect 18580 12960 18670 13200
rect 18910 12960 19000 13200
rect 19240 12960 19330 13200
rect 19570 12960 19920 13200
rect 7610 12870 19920 12960
rect 7610 12630 7780 12870
rect 8020 12630 8110 12870
rect 8350 12630 8440 12870
rect 8680 12630 8770 12870
rect 9010 12630 9100 12870
rect 9340 12630 9430 12870
rect 9670 12630 9760 12870
rect 10000 12630 10090 12870
rect 10330 12630 10420 12870
rect 10660 12630 10750 12870
rect 10990 12630 11080 12870
rect 11320 12630 11410 12870
rect 11650 12630 11740 12870
rect 11980 12630 12070 12870
rect 12310 12630 12400 12870
rect 12640 12630 12730 12870
rect 12970 12630 13060 12870
rect 13300 12630 13390 12870
rect 13630 12630 13720 12870
rect 13960 12630 14050 12870
rect 14290 12630 14380 12870
rect 14620 12630 14710 12870
rect 14950 12630 15040 12870
rect 15280 12630 15370 12870
rect 15610 12630 15700 12870
rect 15940 12630 16030 12870
rect 16270 12630 16360 12870
rect 16600 12630 16690 12870
rect 16930 12630 17020 12870
rect 17260 12630 17350 12870
rect 17590 12630 17680 12870
rect 17920 12630 18010 12870
rect 18250 12630 18340 12870
rect 18580 12630 18670 12870
rect 18910 12630 19000 12870
rect 19240 12630 19330 12870
rect 19570 12630 19920 12870
rect 7610 12540 19920 12630
rect 7610 12300 7780 12540
rect 8020 12300 8110 12540
rect 8350 12300 8440 12540
rect 8680 12300 8770 12540
rect 9010 12300 9100 12540
rect 9340 12300 9430 12540
rect 9670 12300 9760 12540
rect 10000 12300 10090 12540
rect 10330 12300 10420 12540
rect 10660 12300 10750 12540
rect 10990 12300 11080 12540
rect 11320 12300 11410 12540
rect 11650 12300 11740 12540
rect 11980 12300 12070 12540
rect 12310 12300 12400 12540
rect 12640 12300 12730 12540
rect 12970 12300 13060 12540
rect 13300 12300 13390 12540
rect 13630 12300 13720 12540
rect 13960 12300 14050 12540
rect 14290 12300 14380 12540
rect 14620 12300 14710 12540
rect 14950 12300 15040 12540
rect 15280 12300 15370 12540
rect 15610 12300 15700 12540
rect 15940 12300 16030 12540
rect 16270 12300 16360 12540
rect 16600 12300 16690 12540
rect 16930 12300 17020 12540
rect 17260 12300 17350 12540
rect 17590 12300 17680 12540
rect 17920 12300 18010 12540
rect 18250 12300 18340 12540
rect 18580 12300 18670 12540
rect 18910 12300 19000 12540
rect 19240 12300 19330 12540
rect 19570 12300 19920 12540
rect 7610 12210 19920 12300
rect 7610 11970 7780 12210
rect 8020 11970 8110 12210
rect 8350 11970 8440 12210
rect 8680 11970 8770 12210
rect 9010 11970 9100 12210
rect 9340 11970 9430 12210
rect 9670 11970 9760 12210
rect 10000 11970 10090 12210
rect 10330 11970 10420 12210
rect 10660 11970 10750 12210
rect 10990 11970 11080 12210
rect 11320 11970 11410 12210
rect 11650 11970 11740 12210
rect 11980 11970 12070 12210
rect 12310 11970 12400 12210
rect 12640 11970 12730 12210
rect 12970 11970 13060 12210
rect 13300 11970 13390 12210
rect 13630 11970 13720 12210
rect 13960 11970 14050 12210
rect 14290 11970 14380 12210
rect 14620 11970 14710 12210
rect 14950 11970 15040 12210
rect 15280 11970 15370 12210
rect 15610 11970 15700 12210
rect 15940 11970 16030 12210
rect 16270 11970 16360 12210
rect 16600 11970 16690 12210
rect 16930 11970 17020 12210
rect 17260 11970 17350 12210
rect 17590 11970 17680 12210
rect 17920 11970 18010 12210
rect 18250 11970 18340 12210
rect 18580 11970 18670 12210
rect 18910 11970 19000 12210
rect 19240 11970 19330 12210
rect 19570 11970 19920 12210
rect 7610 11880 19920 11970
rect 7610 11640 7780 11880
rect 8020 11640 8110 11880
rect 8350 11640 8440 11880
rect 8680 11640 8770 11880
rect 9010 11640 9100 11880
rect 9340 11640 9430 11880
rect 9670 11640 9760 11880
rect 10000 11640 10090 11880
rect 10330 11640 10420 11880
rect 10660 11640 10750 11880
rect 10990 11640 11080 11880
rect 11320 11640 11410 11880
rect 11650 11640 11740 11880
rect 11980 11640 12070 11880
rect 12310 11640 12400 11880
rect 12640 11640 12730 11880
rect 12970 11640 13060 11880
rect 13300 11640 13390 11880
rect 13630 11640 13720 11880
rect 13960 11640 14050 11880
rect 14290 11640 14380 11880
rect 14620 11640 14710 11880
rect 14950 11640 15040 11880
rect 15280 11640 15370 11880
rect 15610 11640 15700 11880
rect 15940 11640 16030 11880
rect 16270 11640 16360 11880
rect 16600 11640 16690 11880
rect 16930 11640 17020 11880
rect 17260 11640 17350 11880
rect 17590 11640 17680 11880
rect 17920 11640 18010 11880
rect 18250 11640 18340 11880
rect 18580 11640 18670 11880
rect 18910 11640 19000 11880
rect 19240 11640 19330 11880
rect 19570 11640 19920 11880
rect 7610 11550 19920 11640
rect 7610 11310 7780 11550
rect 8020 11310 8110 11550
rect 8350 11310 8440 11550
rect 8680 11310 8770 11550
rect 9010 11310 9100 11550
rect 9340 11310 9430 11550
rect 9670 11310 9760 11550
rect 10000 11310 10090 11550
rect 10330 11310 10420 11550
rect 10660 11310 10750 11550
rect 10990 11310 11080 11550
rect 11320 11310 11410 11550
rect 11650 11310 11740 11550
rect 11980 11310 12070 11550
rect 12310 11310 12400 11550
rect 12640 11310 12730 11550
rect 12970 11310 13060 11550
rect 13300 11310 13390 11550
rect 13630 11310 13720 11550
rect 13960 11310 14050 11550
rect 14290 11310 14380 11550
rect 14620 11310 14710 11550
rect 14950 11310 15040 11550
rect 15280 11310 15370 11550
rect 15610 11310 15700 11550
rect 15940 11310 16030 11550
rect 16270 11310 16360 11550
rect 16600 11310 16690 11550
rect 16930 11310 17020 11550
rect 17260 11310 17350 11550
rect 17590 11310 17680 11550
rect 17920 11310 18010 11550
rect 18250 11310 18340 11550
rect 18580 11310 18670 11550
rect 18910 11310 19000 11550
rect 19240 11310 19330 11550
rect 19570 11310 19920 11550
rect 7610 11220 19920 11310
rect 7610 10980 7780 11220
rect 8020 10980 8110 11220
rect 8350 10980 8440 11220
rect 8680 10980 8770 11220
rect 9010 10980 9100 11220
rect 9340 10980 9430 11220
rect 9670 10980 9760 11220
rect 10000 10980 10090 11220
rect 10330 10980 10420 11220
rect 10660 10980 10750 11220
rect 10990 10980 11080 11220
rect 11320 10980 11410 11220
rect 11650 10980 11740 11220
rect 11980 10980 12070 11220
rect 12310 10980 12400 11220
rect 12640 10980 12730 11220
rect 12970 10980 13060 11220
rect 13300 10980 13390 11220
rect 13630 10980 13720 11220
rect 13960 10980 14050 11220
rect 14290 10980 14380 11220
rect 14620 10980 14710 11220
rect 14950 10980 15040 11220
rect 15280 10980 15370 11220
rect 15610 10980 15700 11220
rect 15940 10980 16030 11220
rect 16270 10980 16360 11220
rect 16600 10980 16690 11220
rect 16930 10980 17020 11220
rect 17260 10980 17350 11220
rect 17590 10980 17680 11220
rect 17920 10980 18010 11220
rect 18250 10980 18340 11220
rect 18580 10980 18670 11220
rect 18910 10980 19000 11220
rect 19240 10980 19330 11220
rect 19570 10980 19920 11220
rect 7610 10890 19920 10980
rect 7610 10650 7780 10890
rect 8020 10650 8110 10890
rect 8350 10650 8440 10890
rect 8680 10650 8770 10890
rect 9010 10650 9100 10890
rect 9340 10650 9430 10890
rect 9670 10650 9760 10890
rect 10000 10650 10090 10890
rect 10330 10650 10420 10890
rect 10660 10650 10750 10890
rect 10990 10650 11080 10890
rect 11320 10650 11410 10890
rect 11650 10650 11740 10890
rect 11980 10650 12070 10890
rect 12310 10650 12400 10890
rect 12640 10650 12730 10890
rect 12970 10650 13060 10890
rect 13300 10650 13390 10890
rect 13630 10650 13720 10890
rect 13960 10650 14050 10890
rect 14290 10650 14380 10890
rect 14620 10650 14710 10890
rect 14950 10650 15040 10890
rect 15280 10650 15370 10890
rect 15610 10650 15700 10890
rect 15940 10650 16030 10890
rect 16270 10650 16360 10890
rect 16600 10650 16690 10890
rect 16930 10650 17020 10890
rect 17260 10650 17350 10890
rect 17590 10650 17680 10890
rect 17920 10650 18010 10890
rect 18250 10650 18340 10890
rect 18580 10650 18670 10890
rect 18910 10650 19000 10890
rect 19240 10650 19330 10890
rect 19570 10650 19920 10890
rect 7610 10560 19920 10650
rect 7610 10320 7780 10560
rect 8020 10320 8110 10560
rect 8350 10320 8440 10560
rect 8680 10320 8770 10560
rect 9010 10320 9100 10560
rect 9340 10320 9430 10560
rect 9670 10320 9760 10560
rect 10000 10320 10090 10560
rect 10330 10320 10420 10560
rect 10660 10320 10750 10560
rect 10990 10320 11080 10560
rect 11320 10320 11410 10560
rect 11650 10320 11740 10560
rect 11980 10320 12070 10560
rect 12310 10320 12400 10560
rect 12640 10320 12730 10560
rect 12970 10320 13060 10560
rect 13300 10320 13390 10560
rect 13630 10320 13720 10560
rect 13960 10320 14050 10560
rect 14290 10320 14380 10560
rect 14620 10320 14710 10560
rect 14950 10320 15040 10560
rect 15280 10320 15370 10560
rect 15610 10320 15700 10560
rect 15940 10320 16030 10560
rect 16270 10320 16360 10560
rect 16600 10320 16690 10560
rect 16930 10320 17020 10560
rect 17260 10320 17350 10560
rect 17590 10320 17680 10560
rect 17920 10320 18010 10560
rect 18250 10320 18340 10560
rect 18580 10320 18670 10560
rect 18910 10320 19000 10560
rect 19240 10320 19330 10560
rect 19570 10320 19920 10560
rect 7610 10230 19920 10320
rect 7610 9990 7780 10230
rect 8020 9990 8110 10230
rect 8350 9990 8440 10230
rect 8680 9990 8770 10230
rect 9010 9990 9100 10230
rect 9340 9990 9430 10230
rect 9670 9990 9760 10230
rect 10000 9990 10090 10230
rect 10330 9990 10420 10230
rect 10660 9990 10750 10230
rect 10990 9990 11080 10230
rect 11320 9990 11410 10230
rect 11650 9990 11740 10230
rect 11980 9990 12070 10230
rect 12310 9990 12400 10230
rect 12640 9990 12730 10230
rect 12970 9990 13060 10230
rect 13300 9990 13390 10230
rect 13630 9990 13720 10230
rect 13960 9990 14050 10230
rect 14290 9990 14380 10230
rect 14620 9990 14710 10230
rect 14950 9990 15040 10230
rect 15280 9990 15370 10230
rect 15610 9990 15700 10230
rect 15940 9990 16030 10230
rect 16270 9990 16360 10230
rect 16600 9990 16690 10230
rect 16930 9990 17020 10230
rect 17260 9990 17350 10230
rect 17590 9990 17680 10230
rect 17920 9990 18010 10230
rect 18250 9990 18340 10230
rect 18580 9990 18670 10230
rect 18910 9990 19000 10230
rect 19240 9990 19330 10230
rect 19570 9990 19920 10230
rect 7610 9900 19920 9990
rect 7610 9660 7780 9900
rect 8020 9660 8110 9900
rect 8350 9660 8440 9900
rect 8680 9660 8770 9900
rect 9010 9660 9100 9900
rect 9340 9660 9430 9900
rect 9670 9660 9760 9900
rect 10000 9660 10090 9900
rect 10330 9660 10420 9900
rect 10660 9660 10750 9900
rect 10990 9660 11080 9900
rect 11320 9660 11410 9900
rect 11650 9660 11740 9900
rect 11980 9660 12070 9900
rect 12310 9660 12400 9900
rect 12640 9660 12730 9900
rect 12970 9660 13060 9900
rect 13300 9660 13390 9900
rect 13630 9660 13720 9900
rect 13960 9660 14050 9900
rect 14290 9660 14380 9900
rect 14620 9660 14710 9900
rect 14950 9660 15040 9900
rect 15280 9660 15370 9900
rect 15610 9660 15700 9900
rect 15940 9660 16030 9900
rect 16270 9660 16360 9900
rect 16600 9660 16690 9900
rect 16930 9660 17020 9900
rect 17260 9660 17350 9900
rect 17590 9660 17680 9900
rect 17920 9660 18010 9900
rect 18250 9660 18340 9900
rect 18580 9660 18670 9900
rect 18910 9660 19000 9900
rect 19240 9660 19330 9900
rect 19570 9660 19920 9900
rect 7610 9570 19920 9660
rect 7610 9330 7780 9570
rect 8020 9330 8110 9570
rect 8350 9330 8440 9570
rect 8680 9330 8770 9570
rect 9010 9330 9100 9570
rect 9340 9330 9430 9570
rect 9670 9330 9760 9570
rect 10000 9330 10090 9570
rect 10330 9330 10420 9570
rect 10660 9330 10750 9570
rect 10990 9330 11080 9570
rect 11320 9330 11410 9570
rect 11650 9330 11740 9570
rect 11980 9330 12070 9570
rect 12310 9330 12400 9570
rect 12640 9330 12730 9570
rect 12970 9330 13060 9570
rect 13300 9330 13390 9570
rect 13630 9330 13720 9570
rect 13960 9330 14050 9570
rect 14290 9330 14380 9570
rect 14620 9330 14710 9570
rect 14950 9330 15040 9570
rect 15280 9330 15370 9570
rect 15610 9330 15700 9570
rect 15940 9330 16030 9570
rect 16270 9330 16360 9570
rect 16600 9330 16690 9570
rect 16930 9330 17020 9570
rect 17260 9330 17350 9570
rect 17590 9330 17680 9570
rect 17920 9330 18010 9570
rect 18250 9330 18340 9570
rect 18580 9330 18670 9570
rect 18910 9330 19000 9570
rect 19240 9330 19330 9570
rect 19570 9330 19920 9570
rect 7610 9240 19920 9330
rect 7610 9000 7780 9240
rect 8020 9000 8110 9240
rect 8350 9000 8440 9240
rect 8680 9000 8770 9240
rect 9010 9000 9100 9240
rect 9340 9000 9430 9240
rect 9670 9000 9760 9240
rect 10000 9000 10090 9240
rect 10330 9000 10420 9240
rect 10660 9000 10750 9240
rect 10990 9000 11080 9240
rect 11320 9000 11410 9240
rect 11650 9000 11740 9240
rect 11980 9000 12070 9240
rect 12310 9000 12400 9240
rect 12640 9000 12730 9240
rect 12970 9000 13060 9240
rect 13300 9000 13390 9240
rect 13630 9000 13720 9240
rect 13960 9000 14050 9240
rect 14290 9000 14380 9240
rect 14620 9000 14710 9240
rect 14950 9000 15040 9240
rect 15280 9000 15370 9240
rect 15610 9000 15700 9240
rect 15940 9000 16030 9240
rect 16270 9000 16360 9240
rect 16600 9000 16690 9240
rect 16930 9000 17020 9240
rect 17260 9000 17350 9240
rect 17590 9000 17680 9240
rect 17920 9000 18010 9240
rect 18250 9000 18340 9240
rect 18580 9000 18670 9240
rect 18910 9000 19000 9240
rect 19240 9000 19330 9240
rect 19570 9000 19920 9240
rect 7610 8830 19920 9000
rect -5020 8500 7340 8510
rect -5020 8430 -4730 8500
rect -4660 8460 -4640 8500
rect -4570 8460 -4550 8500
rect -4480 8460 -4460 8500
rect -4660 8430 -4650 8460
rect -4390 8430 -4370 8500
rect -4300 8460 -4280 8500
rect -4210 8460 -4190 8500
rect -4120 8460 -4100 8500
rect -4030 8430 -4010 8500
rect -3940 8460 -3920 8500
rect -3850 8460 -3830 8500
rect -3760 8460 -3740 8500
rect -3750 8430 -3740 8460
rect -3670 8460 -3650 8500
rect -3580 8460 -3560 8500
rect -3490 8460 -3470 8500
rect -3670 8430 -3660 8460
rect -3400 8430 -3380 8500
rect -3310 8460 -3290 8500
rect -3220 8460 -3200 8500
rect -3130 8460 -3110 8500
rect -3040 8430 -3020 8500
rect -2950 8460 -2930 8500
rect -2860 8460 -2840 8500
rect -2770 8460 -2750 8500
rect -2760 8430 -2750 8460
rect -2680 8460 -2660 8500
rect -2590 8460 -2570 8500
rect -2500 8460 -2480 8500
rect -2680 8430 -2670 8460
rect -2410 8430 -2390 8500
rect -2320 8460 -2300 8500
rect -2230 8460 -2210 8500
rect -2140 8460 -2120 8500
rect -2050 8430 -2030 8500
rect -1960 8460 -1940 8500
rect -1870 8460 -1850 8500
rect -1780 8460 -1720 8500
rect -1770 8430 -1720 8460
rect -1650 8460 -1630 8500
rect -1560 8460 -1540 8500
rect -1470 8460 -1450 8500
rect -1650 8430 -1640 8460
rect -1380 8430 -1360 8500
rect -1290 8460 -1270 8500
rect -1200 8460 -1180 8500
rect -1110 8460 -1090 8500
rect -1020 8430 -1000 8500
rect -930 8460 -910 8500
rect -840 8460 -820 8500
rect -750 8460 -730 8500
rect -740 8430 -730 8460
rect -660 8460 -640 8500
rect -570 8460 -550 8500
rect -480 8460 -460 8500
rect -660 8430 -650 8460
rect -390 8430 -370 8500
rect -300 8460 -280 8500
rect -210 8460 -190 8500
rect -120 8460 -100 8500
rect -30 8430 -10 8500
rect 60 8460 80 8500
rect 150 8460 170 8500
rect 240 8460 260 8500
rect 250 8430 260 8460
rect 330 8460 350 8500
rect 420 8460 440 8500
rect 510 8460 530 8500
rect 330 8430 340 8460
rect 600 8430 620 8500
rect 690 8460 710 8500
rect 780 8460 800 8500
rect 870 8460 890 8500
rect 960 8430 980 8500
rect 1050 8460 1070 8500
rect 1140 8460 1160 8500
rect 1230 8460 1290 8500
rect 1240 8430 1290 8460
rect 1360 8460 1380 8500
rect 1450 8460 1470 8500
rect 1540 8460 1560 8500
rect 1360 8430 1370 8460
rect 1630 8430 1650 8500
rect 1720 8460 1740 8500
rect 1810 8460 1830 8500
rect 1900 8460 1920 8500
rect 1990 8430 2010 8500
rect 2080 8460 2100 8500
rect 2170 8460 2190 8500
rect 2260 8460 2280 8500
rect 2270 8430 2280 8460
rect 2350 8460 2370 8500
rect 2440 8460 2460 8500
rect 2530 8460 2550 8500
rect 2350 8430 2360 8460
rect 2620 8430 2640 8500
rect 2710 8460 2730 8500
rect 2800 8460 2820 8500
rect 2890 8460 2910 8500
rect 2980 8430 3000 8500
rect 3070 8460 3090 8500
rect 3160 8460 3180 8500
rect 3250 8460 3270 8500
rect 3260 8430 3270 8460
rect 3340 8460 3360 8500
rect 3430 8460 3450 8500
rect 3520 8460 3540 8500
rect 3340 8430 3350 8460
rect 3610 8430 3630 8500
rect 3700 8460 3720 8500
rect 3790 8460 3810 8500
rect 3880 8460 3900 8500
rect 3970 8430 3990 8500
rect 4060 8460 4080 8500
rect 4150 8460 4170 8500
rect 4240 8460 4300 8500
rect 4250 8430 4300 8460
rect 4370 8460 4390 8500
rect 4460 8460 4480 8500
rect 4550 8460 4570 8500
rect 4370 8430 4380 8460
rect 4640 8430 4660 8500
rect 4730 8460 4750 8500
rect 4820 8460 4840 8500
rect 4910 8460 4930 8500
rect 5000 8430 5020 8500
rect 5090 8460 5110 8500
rect 5180 8460 5200 8500
rect 5270 8460 5290 8500
rect 5280 8430 5290 8460
rect 5360 8460 5380 8500
rect 5450 8460 5470 8500
rect 5540 8460 5560 8500
rect 5360 8430 5370 8460
rect 5630 8430 5650 8500
rect 5720 8460 5740 8500
rect 5810 8460 5830 8500
rect 5900 8460 5920 8500
rect 5990 8430 6010 8500
rect 6080 8460 6100 8500
rect 6170 8460 6190 8500
rect 6260 8460 6280 8500
rect 6270 8430 6280 8460
rect 6350 8460 6370 8500
rect 6440 8460 6460 8500
rect 6530 8460 6550 8500
rect 6350 8430 6360 8460
rect 6620 8430 6640 8500
rect 6710 8460 6730 8500
rect 6800 8460 6820 8500
rect 6890 8460 6910 8500
rect 6980 8430 7000 8500
rect 7070 8460 7090 8500
rect 7160 8460 7180 8500
rect 7250 8460 7340 8500
rect -5020 8410 -4650 8430
rect -4410 8410 -4320 8430
rect -4080 8410 -3990 8430
rect -3750 8410 -3660 8430
rect -3420 8410 -3330 8430
rect -3090 8410 -3000 8430
rect -2760 8410 -2670 8430
rect -2430 8410 -2340 8430
rect -2100 8410 -2010 8430
rect -1770 8410 -1640 8430
rect -1400 8410 -1310 8430
rect -1070 8410 -980 8430
rect -740 8410 -650 8430
rect -410 8410 -320 8430
rect -80 8410 10 8430
rect 250 8410 340 8430
rect 580 8410 670 8430
rect 910 8410 1000 8430
rect 1240 8410 1370 8430
rect 1610 8410 1700 8430
rect 1940 8410 2030 8430
rect 2270 8410 2360 8430
rect 2600 8410 2690 8430
rect 2930 8410 3020 8430
rect 3260 8410 3350 8430
rect 3590 8410 3680 8430
rect 3920 8410 4010 8430
rect 4250 8410 4380 8430
rect 4620 8410 4710 8430
rect 4950 8410 5040 8430
rect 5280 8410 5370 8430
rect 5610 8410 5700 8430
rect 5940 8410 6030 8430
rect 6270 8410 6360 8430
rect 6600 8410 6690 8430
rect 6930 8410 7020 8430
rect -5020 8340 -4730 8410
rect -4660 8340 -4650 8410
rect -4390 8340 -4370 8410
rect -4030 8340 -4010 8410
rect -3750 8340 -3740 8410
rect -3670 8340 -3660 8410
rect -3400 8340 -3380 8410
rect -3040 8340 -3020 8410
rect -2760 8340 -2750 8410
rect -2680 8340 -2670 8410
rect -2410 8340 -2390 8410
rect -2050 8340 -2030 8410
rect -1770 8340 -1720 8410
rect -1650 8340 -1640 8410
rect -1380 8340 -1360 8410
rect -1020 8340 -1000 8410
rect -740 8340 -730 8410
rect -660 8340 -650 8410
rect -390 8340 -370 8410
rect -30 8340 -10 8410
rect 250 8340 260 8410
rect 330 8340 340 8410
rect 600 8340 620 8410
rect 960 8340 980 8410
rect 1240 8340 1290 8410
rect 1360 8340 1370 8410
rect 1630 8340 1650 8410
rect 1990 8340 2010 8410
rect 2270 8340 2280 8410
rect 2350 8340 2360 8410
rect 2620 8340 2640 8410
rect 2980 8340 3000 8410
rect 3260 8340 3270 8410
rect 3340 8340 3350 8410
rect 3610 8340 3630 8410
rect 3970 8340 3990 8410
rect 4250 8340 4300 8410
rect 4370 8340 4380 8410
rect 4640 8340 4660 8410
rect 5000 8340 5020 8410
rect 5280 8340 5290 8410
rect 5360 8340 5370 8410
rect 5630 8340 5650 8410
rect 5990 8340 6010 8410
rect 6270 8340 6280 8410
rect 6350 8340 6360 8410
rect 6620 8340 6640 8410
rect 6980 8340 7000 8410
rect -5020 8320 -4650 8340
rect -4410 8320 -4320 8340
rect -4080 8320 -3990 8340
rect -3750 8320 -3660 8340
rect -3420 8320 -3330 8340
rect -3090 8320 -3000 8340
rect -2760 8320 -2670 8340
rect -2430 8320 -2340 8340
rect -2100 8320 -2010 8340
rect -1770 8320 -1640 8340
rect -1400 8320 -1310 8340
rect -1070 8320 -980 8340
rect -740 8320 -650 8340
rect -410 8320 -320 8340
rect -80 8320 10 8340
rect 250 8320 340 8340
rect 580 8320 670 8340
rect 910 8320 1000 8340
rect 1240 8320 1370 8340
rect 1610 8320 1700 8340
rect 1940 8320 2030 8340
rect 2270 8320 2360 8340
rect 2600 8320 2690 8340
rect 2930 8320 3020 8340
rect 3260 8320 3350 8340
rect 3590 8320 3680 8340
rect 3920 8320 4010 8340
rect 4250 8320 4380 8340
rect 4620 8320 4710 8340
rect 4950 8320 5040 8340
rect 5280 8320 5370 8340
rect 5610 8320 5700 8340
rect 5940 8320 6030 8340
rect 6270 8320 6360 8340
rect 6600 8320 6690 8340
rect 6930 8320 7020 8340
rect -5020 8250 -4730 8320
rect -4660 8250 -4650 8320
rect -4390 8250 -4370 8320
rect -4030 8250 -4010 8320
rect -3750 8250 -3740 8320
rect -3670 8250 -3660 8320
rect -3400 8250 -3380 8320
rect -3040 8250 -3020 8320
rect -2760 8250 -2750 8320
rect -2680 8250 -2670 8320
rect -2410 8250 -2390 8320
rect -2050 8250 -2030 8320
rect -1770 8250 -1720 8320
rect -1650 8250 -1640 8320
rect -1380 8250 -1360 8320
rect -1020 8250 -1000 8320
rect -740 8250 -730 8320
rect -660 8250 -650 8320
rect -390 8250 -370 8320
rect -30 8250 -10 8320
rect 250 8250 260 8320
rect 330 8250 340 8320
rect 600 8250 620 8320
rect 960 8250 980 8320
rect 1240 8250 1290 8320
rect 1360 8250 1370 8320
rect 1630 8250 1650 8320
rect 1990 8250 2010 8320
rect 2270 8250 2280 8320
rect 2350 8250 2360 8320
rect 2620 8250 2640 8320
rect 2980 8250 3000 8320
rect 3260 8250 3270 8320
rect 3340 8250 3350 8320
rect 3610 8250 3630 8320
rect 3970 8250 3990 8320
rect 4250 8250 4300 8320
rect 4370 8250 4380 8320
rect 4640 8250 4660 8320
rect 5000 8250 5020 8320
rect 5280 8250 5290 8320
rect 5360 8250 5370 8320
rect 5630 8250 5650 8320
rect 5990 8250 6010 8320
rect 6270 8250 6280 8320
rect 6350 8250 6360 8320
rect 6620 8250 6640 8320
rect 6980 8250 7000 8320
rect -5020 8220 -4650 8250
rect -4410 8220 -4320 8250
rect -4080 8220 -3990 8250
rect -3750 8220 -3660 8250
rect -3420 8220 -3330 8250
rect -3090 8220 -3000 8250
rect -2760 8220 -2670 8250
rect -2430 8220 -2340 8250
rect -2100 8220 -2010 8250
rect -1770 8220 -1640 8250
rect -1400 8220 -1310 8250
rect -1070 8220 -980 8250
rect -740 8220 -650 8250
rect -410 8220 -320 8250
rect -80 8220 10 8250
rect 250 8220 340 8250
rect 580 8220 670 8250
rect 910 8220 1000 8250
rect 1240 8220 1370 8250
rect 1610 8220 1700 8250
rect 1940 8220 2030 8250
rect 2270 8220 2360 8250
rect 2600 8220 2690 8250
rect 2930 8220 3020 8250
rect 3260 8220 3350 8250
rect 3590 8220 3680 8250
rect 3920 8220 4010 8250
rect 4250 8220 4380 8250
rect 4620 8220 4710 8250
rect 4950 8220 5040 8250
rect 5280 8220 5370 8250
rect 5610 8220 5700 8250
rect 5940 8220 6030 8250
rect 6270 8220 6360 8250
rect 6600 8220 6690 8250
rect 6930 8220 7020 8250
rect 7260 8220 7340 8460
rect -5020 8190 7340 8220
rect 7020 7910 7340 8190
rect 7020 7840 7040 7910
rect 7110 7840 7140 7910
rect 7210 7840 7240 7910
rect 7310 7840 7340 7910
rect 7020 7820 7340 7840
rect 7020 7750 7040 7820
rect 7110 7750 7140 7820
rect 7210 7750 7240 7820
rect 7310 7750 7340 7820
rect 7020 7730 7340 7750
rect 7560 8500 19920 8510
rect 7560 8460 7650 8500
rect 7720 8460 7740 8500
rect 7810 8460 7830 8500
rect 7560 8220 7640 8460
rect 7900 8430 7920 8500
rect 7990 8460 8010 8500
rect 8080 8460 8100 8500
rect 8170 8460 8190 8500
rect 8260 8430 8280 8500
rect 8350 8460 8370 8500
rect 8440 8460 8460 8500
rect 8530 8460 8550 8500
rect 8540 8430 8550 8460
rect 8620 8460 8640 8500
rect 8710 8460 8730 8500
rect 8800 8460 8820 8500
rect 8620 8430 8630 8460
rect 8890 8430 8910 8500
rect 8980 8460 9000 8500
rect 9070 8460 9090 8500
rect 9160 8460 9180 8500
rect 9250 8430 9270 8500
rect 9340 8460 9360 8500
rect 9430 8460 9450 8500
rect 9520 8460 9540 8500
rect 9530 8430 9540 8460
rect 9610 8460 9630 8500
rect 9700 8460 9720 8500
rect 9790 8460 9810 8500
rect 9610 8430 9620 8460
rect 9880 8430 9900 8500
rect 9970 8460 9990 8500
rect 10060 8460 10080 8500
rect 10150 8460 10170 8500
rect 10240 8430 10260 8500
rect 10330 8460 10350 8500
rect 10420 8460 10440 8500
rect 10510 8460 10530 8500
rect 10520 8430 10530 8460
rect 10600 8460 10660 8500
rect 10730 8460 10750 8500
rect 10820 8460 10840 8500
rect 10600 8430 10650 8460
rect 10910 8430 10930 8500
rect 11000 8460 11020 8500
rect 11090 8460 11110 8500
rect 11180 8460 11200 8500
rect 11270 8430 11290 8500
rect 11360 8460 11380 8500
rect 11450 8460 11470 8500
rect 11540 8460 11560 8500
rect 11550 8430 11560 8460
rect 11630 8460 11650 8500
rect 11720 8460 11740 8500
rect 11810 8460 11830 8500
rect 11630 8430 11640 8460
rect 11900 8430 11920 8500
rect 11990 8460 12010 8500
rect 12080 8460 12100 8500
rect 12170 8460 12190 8500
rect 12260 8430 12280 8500
rect 12350 8460 12370 8500
rect 12440 8460 12460 8500
rect 12530 8460 12550 8500
rect 12540 8430 12550 8460
rect 12620 8460 12640 8500
rect 12710 8460 12730 8500
rect 12800 8460 12820 8500
rect 12620 8430 12630 8460
rect 12890 8430 12910 8500
rect 12980 8460 13000 8500
rect 13070 8460 13090 8500
rect 13160 8460 13180 8500
rect 13250 8430 13270 8500
rect 13340 8460 13360 8500
rect 13430 8460 13450 8500
rect 13520 8460 13540 8500
rect 13530 8430 13540 8460
rect 13610 8460 13670 8500
rect 13740 8460 13760 8500
rect 13830 8460 13850 8500
rect 13610 8430 13660 8460
rect 13920 8430 13940 8500
rect 14010 8460 14030 8500
rect 14100 8460 14120 8500
rect 14190 8460 14210 8500
rect 14280 8430 14300 8500
rect 14370 8460 14390 8500
rect 14460 8460 14480 8500
rect 14550 8460 14570 8500
rect 14560 8430 14570 8460
rect 14640 8460 14660 8500
rect 14730 8460 14750 8500
rect 14820 8460 14840 8500
rect 14640 8430 14650 8460
rect 14910 8430 14930 8500
rect 15000 8460 15020 8500
rect 15090 8460 15110 8500
rect 15180 8460 15200 8500
rect 15270 8430 15290 8500
rect 15360 8460 15380 8500
rect 15450 8460 15470 8500
rect 15540 8460 15560 8500
rect 15550 8430 15560 8460
rect 15630 8460 15650 8500
rect 15720 8460 15740 8500
rect 15810 8460 15830 8500
rect 15630 8430 15640 8460
rect 15900 8430 15920 8500
rect 15990 8460 16010 8500
rect 16080 8460 16100 8500
rect 16170 8460 16190 8500
rect 16260 8430 16280 8500
rect 16350 8460 16370 8500
rect 16440 8460 16460 8500
rect 16530 8460 16550 8500
rect 16540 8430 16550 8460
rect 16620 8460 16680 8500
rect 16750 8460 16770 8500
rect 16840 8460 16860 8500
rect 16620 8430 16670 8460
rect 16930 8430 16950 8500
rect 17020 8460 17040 8500
rect 17110 8460 17130 8500
rect 17200 8460 17220 8500
rect 17290 8430 17310 8500
rect 17380 8460 17400 8500
rect 17470 8460 17490 8500
rect 17560 8460 17580 8500
rect 17570 8430 17580 8460
rect 17650 8460 17670 8500
rect 17740 8460 17760 8500
rect 17830 8460 17850 8500
rect 17650 8430 17660 8460
rect 17920 8430 17940 8500
rect 18010 8460 18030 8500
rect 18100 8460 18120 8500
rect 18190 8460 18210 8500
rect 18280 8430 18300 8500
rect 18370 8460 18390 8500
rect 18460 8460 18480 8500
rect 18550 8460 18570 8500
rect 18560 8430 18570 8460
rect 18640 8460 18660 8500
rect 18730 8460 18750 8500
rect 18820 8460 18840 8500
rect 18640 8430 18650 8460
rect 18910 8430 18930 8500
rect 19000 8460 19020 8500
rect 19090 8460 19110 8500
rect 19180 8460 19200 8500
rect 19270 8430 19290 8500
rect 19360 8460 19380 8500
rect 19450 8460 19470 8500
rect 19540 8460 19560 8500
rect 19550 8430 19560 8460
rect 19630 8430 19920 8500
rect 7880 8410 7970 8430
rect 8210 8410 8300 8430
rect 8540 8410 8630 8430
rect 8870 8410 8960 8430
rect 9200 8410 9290 8430
rect 9530 8410 9620 8430
rect 9860 8410 9950 8430
rect 10190 8410 10280 8430
rect 10520 8410 10650 8430
rect 10890 8410 10980 8430
rect 11220 8410 11310 8430
rect 11550 8410 11640 8430
rect 11880 8410 11970 8430
rect 12210 8410 12300 8430
rect 12540 8410 12630 8430
rect 12870 8410 12960 8430
rect 13200 8410 13290 8430
rect 13530 8410 13660 8430
rect 13900 8410 13990 8430
rect 14230 8410 14320 8430
rect 14560 8410 14650 8430
rect 14890 8410 14980 8430
rect 15220 8410 15310 8430
rect 15550 8410 15640 8430
rect 15880 8410 15970 8430
rect 16210 8410 16300 8430
rect 16540 8410 16670 8430
rect 16910 8410 17000 8430
rect 17240 8410 17330 8430
rect 17570 8410 17660 8430
rect 17900 8410 17990 8430
rect 18230 8410 18320 8430
rect 18560 8410 18650 8430
rect 18890 8410 18980 8430
rect 19220 8410 19310 8430
rect 19550 8410 19920 8430
rect 7900 8340 7920 8410
rect 8260 8340 8280 8410
rect 8540 8340 8550 8410
rect 8620 8340 8630 8410
rect 8890 8340 8910 8410
rect 9250 8340 9270 8410
rect 9530 8340 9540 8410
rect 9610 8340 9620 8410
rect 9880 8340 9900 8410
rect 10240 8340 10260 8410
rect 10520 8340 10530 8410
rect 10600 8340 10650 8410
rect 10910 8340 10930 8410
rect 11270 8340 11290 8410
rect 11550 8340 11560 8410
rect 11630 8340 11640 8410
rect 11900 8340 11920 8410
rect 12260 8340 12280 8410
rect 12540 8340 12550 8410
rect 12620 8340 12630 8410
rect 12890 8340 12910 8410
rect 13250 8340 13270 8410
rect 13530 8340 13540 8410
rect 13610 8340 13660 8410
rect 13920 8340 13940 8410
rect 14280 8340 14300 8410
rect 14560 8340 14570 8410
rect 14640 8340 14650 8410
rect 14910 8340 14930 8410
rect 15270 8340 15290 8410
rect 15550 8340 15560 8410
rect 15630 8340 15640 8410
rect 15900 8340 15920 8410
rect 16260 8340 16280 8410
rect 16540 8340 16550 8410
rect 16620 8340 16670 8410
rect 16930 8340 16950 8410
rect 17290 8340 17310 8410
rect 17570 8340 17580 8410
rect 17650 8340 17660 8410
rect 17920 8340 17940 8410
rect 18280 8340 18300 8410
rect 18560 8340 18570 8410
rect 18640 8340 18650 8410
rect 18910 8340 18930 8410
rect 19270 8340 19290 8410
rect 19550 8340 19560 8410
rect 19630 8340 19920 8410
rect 7880 8320 7970 8340
rect 8210 8320 8300 8340
rect 8540 8320 8630 8340
rect 8870 8320 8960 8340
rect 9200 8320 9290 8340
rect 9530 8320 9620 8340
rect 9860 8320 9950 8340
rect 10190 8320 10280 8340
rect 10520 8320 10650 8340
rect 10890 8320 10980 8340
rect 11220 8320 11310 8340
rect 11550 8320 11640 8340
rect 11880 8320 11970 8340
rect 12210 8320 12300 8340
rect 12540 8320 12630 8340
rect 12870 8320 12960 8340
rect 13200 8320 13290 8340
rect 13530 8320 13660 8340
rect 13900 8320 13990 8340
rect 14230 8320 14320 8340
rect 14560 8320 14650 8340
rect 14890 8320 14980 8340
rect 15220 8320 15310 8340
rect 15550 8320 15640 8340
rect 15880 8320 15970 8340
rect 16210 8320 16300 8340
rect 16540 8320 16670 8340
rect 16910 8320 17000 8340
rect 17240 8320 17330 8340
rect 17570 8320 17660 8340
rect 17900 8320 17990 8340
rect 18230 8320 18320 8340
rect 18560 8320 18650 8340
rect 18890 8320 18980 8340
rect 19220 8320 19310 8340
rect 19550 8320 19920 8340
rect 7900 8250 7920 8320
rect 8260 8250 8280 8320
rect 8540 8250 8550 8320
rect 8620 8250 8630 8320
rect 8890 8250 8910 8320
rect 9250 8250 9270 8320
rect 9530 8250 9540 8320
rect 9610 8250 9620 8320
rect 9880 8250 9900 8320
rect 10240 8250 10260 8320
rect 10520 8250 10530 8320
rect 10600 8250 10650 8320
rect 10910 8250 10930 8320
rect 11270 8250 11290 8320
rect 11550 8250 11560 8320
rect 11630 8250 11640 8320
rect 11900 8250 11920 8320
rect 12260 8250 12280 8320
rect 12540 8250 12550 8320
rect 12620 8250 12630 8320
rect 12890 8250 12910 8320
rect 13250 8250 13270 8320
rect 13530 8250 13540 8320
rect 13610 8250 13660 8320
rect 13920 8250 13940 8320
rect 14280 8250 14300 8320
rect 14560 8250 14570 8320
rect 14640 8250 14650 8320
rect 14910 8250 14930 8320
rect 15270 8250 15290 8320
rect 15550 8250 15560 8320
rect 15630 8250 15640 8320
rect 15900 8250 15920 8320
rect 16260 8250 16280 8320
rect 16540 8250 16550 8320
rect 16620 8250 16670 8320
rect 16930 8250 16950 8320
rect 17290 8250 17310 8320
rect 17570 8250 17580 8320
rect 17650 8250 17660 8320
rect 17920 8250 17940 8320
rect 18280 8250 18300 8320
rect 18560 8250 18570 8320
rect 18640 8250 18650 8320
rect 18910 8250 18930 8320
rect 19270 8250 19290 8320
rect 19550 8250 19560 8320
rect 19630 8250 19920 8320
rect 7880 8220 7970 8250
rect 8210 8220 8300 8250
rect 8540 8220 8630 8250
rect 8870 8220 8960 8250
rect 9200 8220 9290 8250
rect 9530 8220 9620 8250
rect 9860 8220 9950 8250
rect 10190 8220 10280 8250
rect 10520 8220 10650 8250
rect 10890 8220 10980 8250
rect 11220 8220 11310 8250
rect 11550 8220 11640 8250
rect 11880 8220 11970 8250
rect 12210 8220 12300 8250
rect 12540 8220 12630 8250
rect 12870 8220 12960 8250
rect 13200 8220 13290 8250
rect 13530 8220 13660 8250
rect 13900 8220 13990 8250
rect 14230 8220 14320 8250
rect 14560 8220 14650 8250
rect 14890 8220 14980 8250
rect 15220 8220 15310 8250
rect 15550 8220 15640 8250
rect 15880 8220 15970 8250
rect 16210 8220 16300 8250
rect 16540 8220 16670 8250
rect 16910 8220 17000 8250
rect 17240 8220 17330 8250
rect 17570 8220 17660 8250
rect 17900 8220 17990 8250
rect 18230 8220 18320 8250
rect 18560 8220 18650 8250
rect 18890 8220 18980 8250
rect 19220 8220 19310 8250
rect 19550 8220 19920 8250
rect 7560 8190 19920 8220
rect 7560 7910 7880 8190
rect 7560 7840 7590 7910
rect 7660 7840 7690 7910
rect 7760 7840 7790 7910
rect 7860 7840 7880 7910
rect 7560 7820 7880 7840
rect 7560 7750 7590 7820
rect 7660 7750 7690 7820
rect 7760 7750 7790 7820
rect 7860 7750 7880 7820
rect 7560 7730 7880 7750
rect 28700 7830 35460 7910
rect 28700 7590 28780 7830
rect 29020 7590 29110 7830
rect 29350 7590 29440 7830
rect 29680 7590 29770 7830
rect 30010 7590 30100 7830
rect 30340 7590 30430 7830
rect 30670 7590 30760 7830
rect 31000 7590 31090 7830
rect 31330 7590 31420 7830
rect 31660 7590 31750 7830
rect 31990 7590 32080 7830
rect 32320 7590 32410 7830
rect 32650 7590 32740 7830
rect 32980 7590 33070 7830
rect 33310 7590 33400 7830
rect 33640 7590 33730 7830
rect 33970 7590 34060 7830
rect 34300 7590 34390 7830
rect 34630 7590 34720 7830
rect 34960 7590 35050 7830
rect 35290 7590 35460 7830
rect 28700 7500 35460 7590
rect 21060 7270 21540 7290
rect 21060 7210 21110 7270
rect 21480 7210 21540 7270
rect 21060 7140 21090 7210
rect 21490 7140 21540 7210
rect 21060 7100 21110 7140
rect 21480 7100 21540 7140
rect 21060 7030 21090 7100
rect 21490 7030 21540 7100
rect 21060 7000 21540 7030
rect 23460 7270 23940 7290
rect 23460 7210 23510 7270
rect 23880 7210 23940 7270
rect 23460 7140 23490 7210
rect 23890 7140 23940 7210
rect 23460 7100 23510 7140
rect 23880 7100 23940 7140
rect 23460 7030 23490 7100
rect 23890 7030 23940 7100
rect 23460 7000 23940 7030
rect 28700 7260 28780 7500
rect 29020 7260 29110 7500
rect 29350 7260 29440 7500
rect 29680 7260 29770 7500
rect 30010 7260 30100 7500
rect 30340 7260 30430 7500
rect 30670 7260 30760 7500
rect 31000 7260 31090 7500
rect 31330 7260 31420 7500
rect 31660 7260 31750 7500
rect 31990 7260 32080 7500
rect 32320 7260 32410 7500
rect 32650 7260 32740 7500
rect 32980 7260 33070 7500
rect 33310 7260 33400 7500
rect 33640 7260 33730 7500
rect 33970 7260 34060 7500
rect 34300 7260 34390 7500
rect 34630 7260 34720 7500
rect 34960 7260 35050 7500
rect 35290 7260 35460 7500
rect 28700 7170 35460 7260
rect 11760 6940 13360 6960
rect 1540 6910 3140 6930
rect 1540 6850 1720 6910
rect 1960 6850 2050 6910
rect 2290 6850 2390 6910
rect 2630 6850 2720 6910
rect 2960 6850 3140 6910
rect 1540 6780 1570 6850
rect 1640 6780 1680 6850
rect 1970 6780 2010 6850
rect 2300 6780 2340 6850
rect 2630 6780 2670 6850
rect 2960 6780 3000 6850
rect 3070 6780 3140 6850
rect 1540 6740 1720 6780
rect 1960 6740 2050 6780
rect 2290 6740 2390 6780
rect 2630 6740 2720 6780
rect 2960 6740 3140 6780
rect 1540 6670 1570 6740
rect 1640 6670 1680 6740
rect 1970 6670 2010 6740
rect 2300 6670 2340 6740
rect 2630 6670 2670 6740
rect 2960 6670 3000 6740
rect 3070 6670 3140 6740
rect 11760 6880 11940 6940
rect 12180 6880 12270 6940
rect 12510 6880 12610 6940
rect 12850 6880 12940 6940
rect 13180 6880 13360 6940
rect 11760 6810 11790 6880
rect 11860 6810 11900 6880
rect 12190 6810 12230 6880
rect 12520 6810 12560 6880
rect 12850 6810 12890 6880
rect 13180 6810 13220 6880
rect 13290 6810 13360 6880
rect 11760 6770 11940 6810
rect 12180 6770 12270 6810
rect 12510 6770 12610 6810
rect 12850 6770 12940 6810
rect 13180 6770 13360 6810
rect 11760 6700 11790 6770
rect 11860 6700 11900 6770
rect 12190 6700 12230 6770
rect 12520 6700 12560 6770
rect 12850 6700 12890 6770
rect 13180 6700 13220 6770
rect 13290 6700 13360 6770
rect 11760 6670 13360 6700
rect 28700 6930 28780 7170
rect 29020 6930 29110 7170
rect 29350 6930 29440 7170
rect 29680 6930 29770 7170
rect 30010 6930 30100 7170
rect 30340 6930 30430 7170
rect 30670 6930 30760 7170
rect 31000 6930 31090 7170
rect 31330 6930 31420 7170
rect 31660 6930 31750 7170
rect 31990 6930 32080 7170
rect 32320 6930 32410 7170
rect 32650 6930 32740 7170
rect 32980 6930 33070 7170
rect 33310 6930 33400 7170
rect 33640 6930 33730 7170
rect 33970 6930 34060 7170
rect 34300 6930 34390 7170
rect 34630 6930 34720 7170
rect 34960 6930 35050 7170
rect 35290 6930 35460 7170
rect 28700 6840 35460 6930
rect 1540 6640 3140 6670
rect 28700 6600 28780 6840
rect 29020 6600 29110 6840
rect 29350 6600 29440 6840
rect 29680 6600 29770 6840
rect 30010 6600 30100 6840
rect 30340 6600 30430 6840
rect 30670 6600 30760 6840
rect 31000 6600 31090 6840
rect 31330 6600 31420 6840
rect 31660 6600 31750 6840
rect 31990 6600 32080 6840
rect 32320 6600 32410 6840
rect 32650 6600 32740 6840
rect 32980 6600 33070 6840
rect 33310 6600 33400 6840
rect 33640 6600 33730 6840
rect 33970 6600 34060 6840
rect 34300 6600 34390 6840
rect 34630 6600 34720 6840
rect 34960 6600 35050 6840
rect 35290 6600 35460 6840
rect 28700 6510 35460 6600
rect 28700 6320 28780 6510
rect 28320 6300 28780 6320
rect 28320 6230 28340 6300
rect 28410 6230 28450 6300
rect 28520 6270 28780 6300
rect 29020 6270 29110 6510
rect 29350 6270 29440 6510
rect 29680 6270 29770 6510
rect 30010 6270 30100 6510
rect 30340 6270 30430 6510
rect 30670 6270 30760 6510
rect 31000 6270 31090 6510
rect 31330 6270 31420 6510
rect 31660 6270 31750 6510
rect 31990 6270 32080 6510
rect 32320 6270 32410 6510
rect 32650 6270 32740 6510
rect 32980 6270 33070 6510
rect 33310 6270 33400 6510
rect 33640 6270 33730 6510
rect 33970 6270 34060 6510
rect 34300 6270 34390 6510
rect 34630 6270 34720 6510
rect 34960 6270 35050 6510
rect 35290 6270 35460 6510
rect 28520 6230 35460 6270
rect 28320 6180 35460 6230
rect 28320 6170 28780 6180
rect 28320 6100 28340 6170
rect 28410 6100 28450 6170
rect 28520 6100 28780 6170
rect 28320 6040 28780 6100
rect 28320 5970 28340 6040
rect 28410 5970 28450 6040
rect 28520 5970 28780 6040
rect 28320 5950 28780 5970
rect 28700 5940 28780 5950
rect 29020 5940 29110 6180
rect 29350 5940 29440 6180
rect 29680 5940 29770 6180
rect 30010 5940 30100 6180
rect 30340 5940 30430 6180
rect 30670 5940 30760 6180
rect 31000 5940 31090 6180
rect 31330 5940 31420 6180
rect 31660 5940 31750 6180
rect 31990 5940 32080 6180
rect 32320 5940 32410 6180
rect 32650 5940 32740 6180
rect 32980 5940 33070 6180
rect 33310 5940 33400 6180
rect 33640 5940 33730 6180
rect 33970 5940 34060 6180
rect 34300 5940 34390 6180
rect 34630 5940 34720 6180
rect 34960 5940 35050 6180
rect 35290 5940 35460 6180
rect 28700 5850 35460 5940
rect 28700 5610 28780 5850
rect 29020 5610 29110 5850
rect 29350 5610 29440 5850
rect 29680 5610 29770 5850
rect 30010 5610 30100 5850
rect 30340 5610 30430 5850
rect 30670 5610 30760 5850
rect 31000 5610 31090 5850
rect 31330 5610 31420 5850
rect 31660 5610 31750 5850
rect 31990 5610 32080 5850
rect 32320 5610 32410 5850
rect 32650 5610 32740 5850
rect 32980 5610 33070 5850
rect 33310 5610 33400 5850
rect 33640 5610 33730 5850
rect 33970 5610 34060 5850
rect 34300 5610 34390 5850
rect 34630 5610 34720 5850
rect 34960 5610 35050 5850
rect 35290 5610 35460 5850
rect 28700 5520 35460 5610
rect 7400 5390 7490 5410
rect 7400 5320 7410 5390
rect 7480 5320 7490 5390
rect 7400 5280 7490 5320
rect 7400 5210 7410 5280
rect 7480 5210 7490 5280
rect 7400 5185 7490 5210
rect 28700 5280 28780 5520
rect 29020 5280 29110 5520
rect 29350 5280 29440 5520
rect 29680 5280 29770 5520
rect 30010 5280 30100 5520
rect 30340 5280 30430 5520
rect 30670 5280 30760 5520
rect 31000 5280 31090 5520
rect 31330 5280 31420 5520
rect 31660 5280 31750 5520
rect 31990 5280 32080 5520
rect 32320 5280 32410 5520
rect 32650 5280 32740 5520
rect 32980 5280 33070 5520
rect 33310 5280 33400 5520
rect 33640 5280 33730 5520
rect 33970 5280 34060 5520
rect 34300 5280 34390 5520
rect 34630 5280 34720 5520
rect 34960 5280 35050 5520
rect 35290 5280 35460 5520
rect 28700 5190 35460 5280
rect 7400 5170 14790 5185
rect 7400 5100 7410 5170
rect 7480 5100 14790 5170
rect 7400 5075 14790 5100
rect 7400 5060 7490 5075
rect 7400 4990 7410 5060
rect 7480 4990 7490 5060
rect 7400 4950 7490 4990
rect 7400 4880 7410 4950
rect 7480 4880 7490 4950
rect 7400 4860 7490 4880
rect 28700 4950 28780 5190
rect 29020 4950 29110 5190
rect 29350 4950 29440 5190
rect 29680 4950 29770 5190
rect 30010 4950 30100 5190
rect 30340 4950 30430 5190
rect 30670 4950 30760 5190
rect 31000 4950 31090 5190
rect 31330 4950 31420 5190
rect 31660 4950 31750 5190
rect 31990 4950 32080 5190
rect 32320 4950 32410 5190
rect 32650 4950 32740 5190
rect 32980 4950 33070 5190
rect 33310 4950 33400 5190
rect 33640 4950 33730 5190
rect 33970 4950 34060 5190
rect 34300 4950 34390 5190
rect 34630 4950 34720 5190
rect 34960 4950 35050 5190
rect 35290 4950 35460 5190
rect 28700 4860 35460 4950
rect 28700 4620 28780 4860
rect 29020 4620 29110 4860
rect 29350 4620 29440 4860
rect 29680 4620 29770 4860
rect 30010 4620 30100 4860
rect 30340 4620 30430 4860
rect 30670 4620 30760 4860
rect 31000 4620 31090 4860
rect 31330 4620 31420 4860
rect 31660 4620 31750 4860
rect 31990 4620 32080 4860
rect 32320 4620 32410 4860
rect 32650 4620 32740 4860
rect 32980 4620 33070 4860
rect 33310 4620 33400 4860
rect 33640 4620 33730 4860
rect 33970 4620 34060 4860
rect 34300 4620 34390 4860
rect 34630 4620 34720 4860
rect 34960 4620 35050 4860
rect 35290 4620 35460 4860
rect 28700 4530 35460 4620
rect 28700 4290 28780 4530
rect 29020 4290 29110 4530
rect 29350 4290 29440 4530
rect 29680 4290 29770 4530
rect 30010 4290 30100 4530
rect 30340 4290 30430 4530
rect 30670 4290 30760 4530
rect 31000 4290 31090 4530
rect 31330 4290 31420 4530
rect 31660 4290 31750 4530
rect 31990 4290 32080 4530
rect 32320 4290 32410 4530
rect 32650 4290 32740 4530
rect 32980 4290 33070 4530
rect 33310 4290 33400 4530
rect 33640 4290 33730 4530
rect 33970 4290 34060 4530
rect 34300 4290 34390 4530
rect 34630 4290 34720 4530
rect 34960 4290 35050 4530
rect 35290 4290 35460 4530
rect 28700 4200 35460 4290
rect 28700 3960 28780 4200
rect 29020 3960 29110 4200
rect 29350 3960 29440 4200
rect 29680 3960 29770 4200
rect 30010 3960 30100 4200
rect 30340 3960 30430 4200
rect 30670 3960 30760 4200
rect 31000 3960 31090 4200
rect 31330 3960 31420 4200
rect 31660 3960 31750 4200
rect 31990 3960 32080 4200
rect 32320 3960 32410 4200
rect 32650 3960 32740 4200
rect 32980 3960 33070 4200
rect 33310 3960 33400 4200
rect 33640 3960 33730 4200
rect 33970 3960 34060 4200
rect 34300 3960 34390 4200
rect 34630 3960 34720 4200
rect 34960 3960 35050 4200
rect 35290 3960 35460 4200
rect 28700 3870 35460 3960
rect 28700 3630 28780 3870
rect 29020 3630 29110 3870
rect 29350 3630 29440 3870
rect 29680 3630 29770 3870
rect 30010 3630 30100 3870
rect 30340 3630 30430 3870
rect 30670 3630 30760 3870
rect 31000 3630 31090 3870
rect 31330 3630 31420 3870
rect 31660 3630 31750 3870
rect 31990 3630 32080 3870
rect 32320 3630 32410 3870
rect 32650 3630 32740 3870
rect 32980 3630 33070 3870
rect 33310 3630 33400 3870
rect 33640 3630 33730 3870
rect 33970 3630 34060 3870
rect 34300 3630 34390 3870
rect 34630 3630 34720 3870
rect 34960 3630 35050 3870
rect 35290 3630 35460 3870
rect 28700 3540 35460 3630
rect 22300 3360 22630 3380
rect 22300 3290 22320 3360
rect 22390 3290 22430 3360
rect 22500 3290 22540 3360
rect 22610 3290 22630 3360
rect 22300 3250 22630 3290
rect 22300 3236 22320 3250
rect 22284 3180 22320 3236
rect 22390 3180 22430 3250
rect 22500 3180 22540 3250
rect 22610 3236 22630 3250
rect 28700 3300 28780 3540
rect 29020 3300 29110 3540
rect 29350 3300 29440 3540
rect 29680 3300 29770 3540
rect 30010 3300 30100 3540
rect 30340 3300 30430 3540
rect 30670 3300 30760 3540
rect 31000 3300 31090 3540
rect 31330 3300 31420 3540
rect 31660 3300 31750 3540
rect 31990 3300 32080 3540
rect 32320 3300 32410 3540
rect 32650 3300 32740 3540
rect 32980 3300 33070 3540
rect 33310 3300 33400 3540
rect 33640 3300 33730 3540
rect 33970 3300 34060 3540
rect 34300 3300 34390 3540
rect 34630 3300 34720 3540
rect 34960 3300 35050 3540
rect 35290 3300 35460 3540
rect 22610 3180 28077 3236
rect 22284 3140 28077 3180
rect 22284 3103 22320 3140
rect 22300 3070 22320 3103
rect 22390 3070 22430 3140
rect 22500 3070 22540 3140
rect 22610 3103 28077 3140
rect 22610 3070 22630 3103
rect 22300 3050 22630 3070
rect 20020 2600 20500 2630
rect 20020 2530 20070 2600
rect 20470 2530 20500 2600
rect 20020 2490 20080 2530
rect 20450 2490 20500 2530
rect 20020 2420 20070 2490
rect 20470 2420 20500 2490
rect 20020 2360 20080 2420
rect 20450 2360 20500 2420
rect 20020 2340 20500 2360
rect 24500 2600 24980 2630
rect 24500 2530 24550 2600
rect 24950 2530 24980 2600
rect 24500 2490 24560 2530
rect 24930 2490 24980 2530
rect 24500 2420 24550 2490
rect 24950 2420 24980 2490
rect 24500 2360 24560 2420
rect 24930 2360 24980 2420
rect 24500 2340 24980 2360
rect 14590 1160 15150 1180
rect 14590 1090 14600 1160
rect 14670 1090 14700 1160
rect 14770 1090 14810 1160
rect 14880 1090 15150 1160
rect 14590 1050 16685 1090
rect 14590 980 14600 1050
rect 14670 980 14700 1050
rect 14770 980 14810 1050
rect 14880 980 16685 1050
rect 14590 960 16685 980
rect 14590 940 15150 960
rect 14590 870 14600 940
rect 14670 870 14700 940
rect 14770 870 14810 940
rect 14880 870 15150 940
rect 14590 850 15150 870
rect 1080 -790 2680 -760
rect 1080 -860 1150 -790
rect 1220 -860 1260 -790
rect 1550 -860 1590 -790
rect 1880 -860 1920 -790
rect 2210 -860 2250 -790
rect 2540 -860 2580 -790
rect 2650 -860 2680 -790
rect 1080 -900 1260 -860
rect 1500 -900 1590 -860
rect 1830 -900 1930 -860
rect 2170 -900 2260 -860
rect 2500 -900 2680 -860
rect 1080 -970 1150 -900
rect 1220 -970 1260 -900
rect 1550 -970 1590 -900
rect 1880 -970 1920 -900
rect 2210 -970 2250 -900
rect 2540 -970 2580 -900
rect 2650 -970 2680 -900
rect 1080 -1030 1260 -970
rect 1500 -1030 1590 -970
rect 1830 -1030 1930 -970
rect 2170 -1030 2260 -970
rect 2500 -1030 2680 -970
rect 1080 -1050 2680 -1030
rect 12220 -790 13820 -760
rect 12220 -860 12250 -790
rect 12320 -860 12360 -790
rect 12650 -860 12690 -790
rect 12980 -860 13020 -790
rect 13310 -860 13350 -790
rect 13640 -860 13680 -790
rect 13750 -860 13820 -790
rect 12220 -900 12400 -860
rect 12640 -900 12730 -860
rect 12970 -900 13070 -860
rect 13310 -900 13400 -860
rect 13640 -900 13820 -860
rect 12220 -970 12250 -900
rect 12320 -970 12360 -900
rect 12650 -970 12690 -900
rect 12980 -970 13020 -900
rect 13310 -970 13350 -900
rect 13640 -970 13680 -900
rect 13750 -970 13820 -900
rect 12220 -1030 12400 -970
rect 12640 -1030 12730 -970
rect 12970 -1030 13070 -970
rect 13310 -1030 13400 -970
rect 13640 -1030 13820 -970
rect 12220 -1050 13820 -1030
rect 1540 -2720 3140 -2700
rect 1540 -2780 1720 -2720
rect 1960 -2780 2050 -2720
rect 2290 -2780 2390 -2720
rect 2630 -2780 2720 -2720
rect 2960 -2780 3140 -2720
rect 1540 -2850 1570 -2780
rect 1640 -2850 1680 -2780
rect 1970 -2850 2010 -2780
rect 2300 -2850 2340 -2780
rect 2630 -2850 2670 -2780
rect 2960 -2850 3000 -2780
rect 3070 -2850 3140 -2780
rect 1540 -2890 1720 -2850
rect 1960 -2890 2050 -2850
rect 2290 -2890 2390 -2850
rect 2630 -2890 2720 -2850
rect 2960 -2890 3140 -2850
rect 1540 -2960 1570 -2890
rect 1640 -2960 1680 -2890
rect 1970 -2960 2010 -2890
rect 2300 -2960 2340 -2890
rect 2630 -2960 2670 -2890
rect 2960 -2960 3000 -2890
rect 3070 -2960 3140 -2890
rect 1540 -2990 3140 -2960
rect 11760 -2720 13360 -2700
rect 11760 -2780 11940 -2720
rect 12180 -2780 12270 -2720
rect 12510 -2780 12610 -2720
rect 12850 -2780 12940 -2720
rect 13180 -2780 13360 -2720
rect 11760 -2850 11790 -2780
rect 11860 -2850 11900 -2780
rect 12190 -2850 12230 -2780
rect 12520 -2850 12560 -2780
rect 12850 -2850 12890 -2780
rect 13180 -2850 13220 -2780
rect 13290 -2850 13360 -2780
rect 11760 -2890 11940 -2850
rect 12180 -2890 12270 -2850
rect 12510 -2890 12610 -2850
rect 12850 -2890 12940 -2850
rect 13180 -2890 13360 -2850
rect 11760 -2960 11790 -2890
rect 11860 -2960 11900 -2890
rect 12190 -2960 12230 -2890
rect 12520 -2960 12560 -2890
rect 12850 -2960 12890 -2890
rect 13180 -2960 13220 -2890
rect 13290 -2960 13360 -2890
rect 11760 -2990 13360 -2960
rect -1860 -4260 -250 -4050
rect -1860 -4500 -1650 -4260
rect -1410 -4500 -1320 -4260
rect -1080 -4500 -990 -4260
rect -750 -4500 -660 -4260
rect -420 -4500 -250 -4260
rect -1860 -4590 -250 -4500
rect -1860 -4830 -1650 -4590
rect -1410 -4830 -1320 -4590
rect -1080 -4830 -990 -4590
rect -750 -4830 -660 -4590
rect -420 -4830 -250 -4590
rect -1860 -4920 -250 -4830
rect -1860 -5160 -1650 -4920
rect -1410 -5160 -1320 -4920
rect -1080 -5160 -990 -4920
rect -750 -5160 -660 -4920
rect -420 -5160 -250 -4920
rect -1860 -5180 -250 -5160
rect -2220 -5240 -250 -5180
rect -2220 -5310 -2140 -5240
rect -2070 -5310 -2030 -5240
rect -1960 -5250 -250 -5240
rect -1960 -5310 -1650 -5250
rect -2220 -5350 -1650 -5310
rect -2220 -5420 -2140 -5350
rect -2070 -5420 -2030 -5350
rect -1960 -5420 -1650 -5350
rect -2220 -5460 -1650 -5420
rect -2220 -5530 -2140 -5460
rect -2070 -5530 -2030 -5460
rect -1960 -5490 -1650 -5460
rect -1410 -5490 -1320 -5250
rect -1080 -5490 -990 -5250
rect -750 -5490 -660 -5250
rect -420 -5490 -250 -5250
rect -1960 -5530 -250 -5490
rect -170 -4230 150 -4220
rect -170 -4300 -160 -4230
rect -90 -4250 -70 -4230
rect 0 -4250 20 -4230
rect 90 -4250 150 -4230
rect -170 -4320 -120 -4300
rect -170 -4390 -160 -4320
rect -170 -4410 -120 -4390
rect -170 -4480 -160 -4410
rect -170 -4490 -120 -4480
rect 120 -4490 150 -4250
rect -170 -4500 150 -4490
rect -170 -4570 -160 -4500
rect -90 -4570 -70 -4500
rect 0 -4570 20 -4500
rect 90 -4570 150 -4500
rect -170 -4580 150 -4570
rect -170 -4590 -120 -4580
rect -170 -4660 -160 -4590
rect -170 -4680 -120 -4660
rect -170 -4750 -160 -4680
rect -170 -4770 -120 -4750
rect -170 -4840 -160 -4770
rect 120 -4820 150 -4580
rect -90 -4840 -70 -4820
rect 0 -4840 20 -4820
rect 90 -4840 150 -4820
rect -170 -4860 150 -4840
rect -170 -4930 -160 -4860
rect -90 -4910 -70 -4860
rect 0 -4910 20 -4860
rect 90 -4910 150 -4860
rect 7290 -4560 7620 -4540
rect 7290 -4630 7310 -4560
rect 7380 -4630 7420 -4560
rect 7490 -4630 7530 -4560
rect 7600 -4600 7620 -4560
rect 7600 -4630 15780 -4600
rect 7290 -4670 15780 -4630
rect 7290 -4740 7310 -4670
rect 7380 -4740 7420 -4670
rect 7490 -4740 7530 -4670
rect 7600 -4740 15780 -4670
rect 7290 -4760 15780 -4740
rect 7290 -4780 7620 -4760
rect 7290 -4850 7310 -4780
rect 7380 -4850 7420 -4780
rect 7490 -4850 7530 -4780
rect 7600 -4850 7620 -4780
rect 7290 -4870 7620 -4850
rect -170 -4950 -120 -4930
rect -170 -5020 -160 -4950
rect -170 -5040 -120 -5020
rect -170 -5110 -160 -5040
rect -170 -5130 -120 -5110
rect -170 -5200 -160 -5130
rect 120 -5150 150 -4910
rect -90 -5200 -70 -5150
rect 0 -5200 20 -5150
rect 90 -5200 150 -5150
rect -170 -5220 150 -5200
rect -170 -5290 -160 -5220
rect -90 -5240 -70 -5220
rect 0 -5240 20 -5220
rect 90 -5240 150 -5220
rect -170 -5310 -120 -5290
rect -170 -5380 -160 -5310
rect -170 -5400 -120 -5380
rect -170 -5470 -160 -5400
rect -170 -5480 -120 -5470
rect 120 -5480 150 -5240
rect -170 -5510 150 -5480
rect -2220 -5570 -250 -5530
rect -2220 -5640 -2140 -5570
rect -2070 -5640 -2030 -5570
rect -1960 -5640 -250 -5570
rect -2220 -5660 -250 -5640
rect 16575 -5915 16685 960
rect 21060 980 21540 1000
rect 21060 920 21110 980
rect 21480 920 21540 980
rect 21060 850 21090 920
rect 21490 850 21540 920
rect 21060 810 21110 850
rect 21480 810 21540 850
rect 21060 740 21090 810
rect 21490 740 21540 810
rect 21060 710 21540 740
rect 23460 980 23940 1000
rect 23460 920 23510 980
rect 23880 920 23940 980
rect 23460 850 23490 920
rect 23890 850 23940 920
rect 23460 810 23510 850
rect 23880 810 23940 850
rect 23460 740 23490 810
rect 23890 740 23940 810
rect 23460 710 23940 740
rect 22320 -3050 22650 -3030
rect 22320 -3120 22340 -3050
rect 22410 -3120 22450 -3050
rect 22520 -3120 22560 -3050
rect 22630 -3120 22650 -3050
rect 22320 -3125 22650 -3120
rect 27944 -3125 28077 3103
rect 28700 3210 35460 3300
rect 28700 2970 28780 3210
rect 29020 2970 29110 3210
rect 29350 2970 29440 3210
rect 29680 2970 29770 3210
rect 30010 2970 30100 3210
rect 30340 2970 30430 3210
rect 30670 2970 30760 3210
rect 31000 2970 31090 3210
rect 31330 2970 31420 3210
rect 31660 2970 31750 3210
rect 31990 2970 32080 3210
rect 32320 2970 32410 3210
rect 32650 2970 32740 3210
rect 32980 2970 33070 3210
rect 33310 2970 33400 3210
rect 33640 2970 33730 3210
rect 33970 2970 34060 3210
rect 34300 2970 34390 3210
rect 34630 2970 34720 3210
rect 34960 2970 35050 3210
rect 35290 2970 35460 3210
rect 28700 2880 35460 2970
rect 28700 2640 28780 2880
rect 29020 2640 29110 2880
rect 29350 2640 29440 2880
rect 29680 2640 29770 2880
rect 30010 2640 30100 2880
rect 30340 2640 30430 2880
rect 30670 2640 30760 2880
rect 31000 2640 31090 2880
rect 31330 2640 31420 2880
rect 31660 2640 31750 2880
rect 31990 2640 32080 2880
rect 32320 2640 32410 2880
rect 32650 2640 32740 2880
rect 32980 2640 33070 2880
rect 33310 2640 33400 2880
rect 33640 2640 33730 2880
rect 33970 2640 34060 2880
rect 34300 2640 34390 2880
rect 34630 2640 34720 2880
rect 34960 2640 35050 2880
rect 35290 2640 35460 2880
rect 28700 2550 35460 2640
rect 28700 2310 28780 2550
rect 29020 2310 29110 2550
rect 29350 2310 29440 2550
rect 29680 2310 29770 2550
rect 30010 2310 30100 2550
rect 30340 2310 30430 2550
rect 30670 2310 30760 2550
rect 31000 2310 31090 2550
rect 31330 2310 31420 2550
rect 31660 2310 31750 2550
rect 31990 2310 32080 2550
rect 32320 2310 32410 2550
rect 32650 2310 32740 2550
rect 32980 2310 33070 2550
rect 33310 2310 33400 2550
rect 33640 2310 33730 2550
rect 33970 2310 34060 2550
rect 34300 2310 34390 2550
rect 34630 2310 34720 2550
rect 34960 2310 35050 2550
rect 35290 2310 35460 2550
rect 28700 2220 35460 2310
rect 28700 1980 28780 2220
rect 29020 1980 29110 2220
rect 29350 1980 29440 2220
rect 29680 1980 29770 2220
rect 30010 1980 30100 2220
rect 30340 1980 30430 2220
rect 30670 1980 30760 2220
rect 31000 1980 31090 2220
rect 31330 1980 31420 2220
rect 31660 1980 31750 2220
rect 31990 1980 32080 2220
rect 32320 1980 32410 2220
rect 32650 1980 32740 2220
rect 32980 1980 33070 2220
rect 33310 1980 33400 2220
rect 33640 1980 33730 2220
rect 33970 1980 34060 2220
rect 34300 1980 34390 2220
rect 34630 1980 34720 2220
rect 34960 1980 35050 2220
rect 35290 1980 35460 2220
rect 28700 1890 35460 1980
rect 28700 1650 28780 1890
rect 29020 1650 29110 1890
rect 29350 1650 29440 1890
rect 29680 1650 29770 1890
rect 30010 1650 30100 1890
rect 30340 1650 30430 1890
rect 30670 1650 30760 1890
rect 31000 1650 31090 1890
rect 31330 1650 31420 1890
rect 31660 1650 31750 1890
rect 31990 1650 32080 1890
rect 32320 1650 32410 1890
rect 32650 1650 32740 1890
rect 32980 1650 33070 1890
rect 33310 1650 33400 1890
rect 33640 1650 33730 1890
rect 33970 1650 34060 1890
rect 34300 1650 34390 1890
rect 34630 1650 34720 1890
rect 34960 1650 35050 1890
rect 35290 1650 35460 1890
rect 28700 1560 35460 1650
rect 28700 1320 28780 1560
rect 29020 1320 29110 1560
rect 29350 1320 29440 1560
rect 29680 1320 29770 1560
rect 30010 1320 30100 1560
rect 30340 1320 30430 1560
rect 30670 1320 30760 1560
rect 31000 1320 31090 1560
rect 31330 1320 31420 1560
rect 31660 1320 31750 1560
rect 31990 1320 32080 1560
rect 32320 1320 32410 1560
rect 32650 1320 32740 1560
rect 32980 1320 33070 1560
rect 33310 1320 33400 1560
rect 33640 1320 33730 1560
rect 33970 1320 34060 1560
rect 34300 1320 34390 1560
rect 34630 1320 34720 1560
rect 34960 1320 35050 1560
rect 35290 1320 35460 1560
rect 28700 1150 35460 1320
rect 35780 7820 36100 7910
rect 35780 7750 35790 7820
rect 35860 7770 35880 7820
rect 35950 7770 35970 7820
rect 36040 7770 36100 7820
rect 35780 7730 35830 7750
rect 35780 7660 35790 7730
rect 35780 7640 35830 7660
rect 35780 7570 35790 7640
rect 35780 7550 35830 7570
rect 35780 7480 35790 7550
rect 36070 7530 36100 7770
rect 35860 7480 35880 7530
rect 35950 7480 35970 7530
rect 36040 7480 36100 7530
rect 35780 7460 36100 7480
rect 35780 7390 35790 7460
rect 35860 7440 35880 7460
rect 35950 7440 35970 7460
rect 36040 7440 36100 7460
rect 35780 7370 35830 7390
rect 35780 7300 35790 7370
rect 35780 7280 35830 7300
rect 35780 7210 35790 7280
rect 35780 7200 35830 7210
rect 36070 7200 36100 7440
rect 35780 7150 36100 7200
rect 35780 7080 35790 7150
rect 35860 7080 35880 7150
rect 35950 7080 35970 7150
rect 36040 7080 36100 7150
rect 35780 7070 36100 7080
rect 35780 7060 35830 7070
rect 35780 6990 35790 7060
rect 35780 6970 35830 6990
rect 35780 6900 35790 6970
rect 35780 6880 35830 6900
rect 35780 6810 35790 6880
rect 36070 6830 36100 7070
rect 35860 6810 35880 6830
rect 35950 6810 35970 6830
rect 36040 6810 36100 6830
rect 35780 6790 36100 6810
rect 35780 6720 35790 6790
rect 35860 6740 35880 6790
rect 35950 6740 35970 6790
rect 36040 6740 36100 6790
rect 35780 6700 35830 6720
rect 35780 6630 35790 6700
rect 35780 6610 35830 6630
rect 35780 6540 35790 6610
rect 35780 6520 35830 6540
rect 35780 6450 35790 6520
rect 36070 6500 36100 6740
rect 35860 6450 35880 6500
rect 35950 6450 35970 6500
rect 36040 6450 36100 6500
rect 35780 6430 36100 6450
rect 35780 6360 35790 6430
rect 35860 6410 35880 6430
rect 35950 6410 35970 6430
rect 36040 6410 36100 6430
rect 35780 6340 35830 6360
rect 35780 6270 35790 6340
rect 35780 6250 35830 6270
rect 35780 6180 35790 6250
rect 35780 6170 35830 6180
rect 36070 6170 36100 6410
rect 35780 6160 36100 6170
rect 35780 6090 35790 6160
rect 35860 6090 35880 6160
rect 35950 6090 35970 6160
rect 36040 6090 36100 6160
rect 35780 6080 36100 6090
rect 35780 6070 35830 6080
rect 35780 6000 35790 6070
rect 35780 5980 35830 6000
rect 35780 5910 35790 5980
rect 35780 5890 35830 5910
rect 35780 5820 35790 5890
rect 36070 5840 36100 6080
rect 35860 5820 35880 5840
rect 35950 5820 35970 5840
rect 36040 5820 36100 5840
rect 35780 5800 36100 5820
rect 35780 5730 35790 5800
rect 35860 5750 35880 5800
rect 35950 5750 35970 5800
rect 36040 5750 36100 5800
rect 35780 5710 35830 5730
rect 35780 5640 35790 5710
rect 35780 5620 35830 5640
rect 35780 5550 35790 5620
rect 35780 5530 35830 5550
rect 35780 5460 35790 5530
rect 36070 5510 36100 5750
rect 35860 5460 35880 5510
rect 35950 5460 35970 5510
rect 36040 5460 36100 5510
rect 35780 5440 36100 5460
rect 35780 5370 35790 5440
rect 35860 5420 35880 5440
rect 35950 5420 35970 5440
rect 36040 5420 36100 5440
rect 35780 5350 35830 5370
rect 35780 5280 35790 5350
rect 35780 5260 35830 5280
rect 35780 5190 35790 5260
rect 35780 5180 35830 5190
rect 36070 5180 36100 5420
rect 35780 5170 36100 5180
rect 35780 5100 35790 5170
rect 35860 5100 35880 5170
rect 35950 5100 35970 5170
rect 36040 5100 36100 5170
rect 35780 5090 36100 5100
rect 35780 5080 35830 5090
rect 35780 5010 35790 5080
rect 35780 4990 35830 5010
rect 35780 4920 35790 4990
rect 35780 4900 35830 4920
rect 35780 4830 35790 4900
rect 36070 4850 36100 5090
rect 35860 4830 35880 4850
rect 35950 4830 35970 4850
rect 36040 4830 36100 4850
rect 35780 4810 36100 4830
rect 35780 4740 35790 4810
rect 35860 4760 35880 4810
rect 35950 4760 35970 4810
rect 36040 4760 36100 4810
rect 35780 4720 35830 4740
rect 35780 4650 35790 4720
rect 35780 4630 35830 4650
rect 35780 4560 35790 4630
rect 35780 4540 35830 4560
rect 35780 4470 35790 4540
rect 36070 4520 36100 4760
rect 35860 4470 35880 4520
rect 35950 4470 35970 4520
rect 36040 4470 36100 4520
rect 35780 4450 36100 4470
rect 35780 4380 35790 4450
rect 35860 4430 35880 4450
rect 35950 4430 35970 4450
rect 36040 4430 36100 4450
rect 35780 4360 35830 4380
rect 35780 4290 35790 4360
rect 35780 4270 35830 4290
rect 35780 4200 35790 4270
rect 35780 4190 35830 4200
rect 36070 4190 36100 4430
rect 35780 4140 36100 4190
rect 35780 4070 35790 4140
rect 35860 4070 35880 4140
rect 35950 4070 35970 4140
rect 36040 4070 36100 4140
rect 35780 4060 36100 4070
rect 35780 4050 35830 4060
rect 35780 3980 35790 4050
rect 35780 3960 35830 3980
rect 35780 3890 35790 3960
rect 35780 3870 35830 3890
rect 35780 3800 35790 3870
rect 36070 3820 36100 4060
rect 35860 3800 35880 3820
rect 35950 3800 35970 3820
rect 36040 3800 36100 3820
rect 35780 3780 36100 3800
rect 35780 3710 35790 3780
rect 35860 3730 35880 3780
rect 35950 3730 35970 3780
rect 36040 3730 36100 3780
rect 35780 3690 35830 3710
rect 35780 3620 35790 3690
rect 35780 3600 35830 3620
rect 35780 3530 35790 3600
rect 35780 3510 35830 3530
rect 35780 3440 35790 3510
rect 36070 3490 36100 3730
rect 35860 3440 35880 3490
rect 35950 3440 35970 3490
rect 36040 3440 36100 3490
rect 35780 3420 36100 3440
rect 35780 3350 35790 3420
rect 35860 3400 35880 3420
rect 35950 3400 35970 3420
rect 36040 3400 36100 3420
rect 35780 3330 35830 3350
rect 35780 3260 35790 3330
rect 35780 3240 35830 3260
rect 35780 3170 35790 3240
rect 35780 3160 35830 3170
rect 36070 3160 36100 3400
rect 35780 3150 36100 3160
rect 35780 3080 35790 3150
rect 35860 3080 35880 3150
rect 35950 3080 35970 3150
rect 36040 3080 36100 3150
rect 35780 3070 36100 3080
rect 35780 3060 35830 3070
rect 35780 2990 35790 3060
rect 35780 2970 35830 2990
rect 35780 2900 35790 2970
rect 35780 2880 35830 2900
rect 35780 2810 35790 2880
rect 36070 2830 36100 3070
rect 35860 2810 35880 2830
rect 35950 2810 35970 2830
rect 36040 2810 36100 2830
rect 35780 2790 36100 2810
rect 35780 2720 35790 2790
rect 35860 2740 35880 2790
rect 35950 2740 35970 2790
rect 36040 2740 36100 2790
rect 35780 2700 35830 2720
rect 35780 2630 35790 2700
rect 35780 2610 35830 2630
rect 35780 2540 35790 2610
rect 35780 2520 35830 2540
rect 35780 2450 35790 2520
rect 36070 2500 36100 2740
rect 35860 2450 35880 2500
rect 35950 2450 35970 2500
rect 36040 2450 36100 2500
rect 35780 2430 36100 2450
rect 35780 2360 35790 2430
rect 35860 2410 35880 2430
rect 35950 2410 35970 2430
rect 36040 2410 36100 2430
rect 35780 2340 35830 2360
rect 35780 2270 35790 2340
rect 35780 2250 35830 2270
rect 35780 2180 35790 2250
rect 35780 2170 35830 2180
rect 36070 2170 36100 2410
rect 35780 2160 36100 2170
rect 35780 2090 35790 2160
rect 35860 2090 35880 2160
rect 35950 2090 35970 2160
rect 36040 2090 36100 2160
rect 35780 2080 36100 2090
rect 35780 2070 35830 2080
rect 35780 2000 35790 2070
rect 35780 1980 35830 2000
rect 35780 1910 35790 1980
rect 35780 1890 35830 1910
rect 35780 1820 35790 1890
rect 36070 1840 36100 2080
rect 35860 1820 35880 1840
rect 35950 1820 35970 1840
rect 36040 1820 36100 1840
rect 35780 1800 36100 1820
rect 35780 1730 35790 1800
rect 35860 1750 35880 1800
rect 35950 1750 35970 1800
rect 36040 1750 36100 1800
rect 35780 1710 35830 1730
rect 35780 1640 35790 1710
rect 35780 1620 35830 1640
rect 35780 1550 35790 1620
rect 35780 1530 35830 1550
rect 35780 1460 35790 1530
rect 36070 1510 36100 1750
rect 35860 1460 35880 1510
rect 35950 1460 35970 1510
rect 36040 1460 36100 1510
rect 35780 1440 36100 1460
rect 35780 1370 35790 1440
rect 35860 1420 35880 1440
rect 35950 1420 35970 1440
rect 36040 1420 36100 1440
rect 35780 1350 35830 1370
rect 35780 1280 35790 1350
rect 35780 1260 35830 1280
rect 35780 1190 35790 1260
rect 35780 1180 35830 1190
rect 36070 1180 36100 1420
rect 35780 1150 36100 1180
rect 28700 230 35460 310
rect 28700 20 28780 230
rect 28320 0 28780 20
rect 28320 -70 28340 0
rect 28410 -70 28450 0
rect 28520 -10 28780 0
rect 29020 -10 29110 230
rect 29350 -10 29440 230
rect 29680 -10 29770 230
rect 30010 -10 30100 230
rect 30340 -10 30430 230
rect 30670 -10 30760 230
rect 31000 -10 31090 230
rect 31330 -10 31420 230
rect 31660 -10 31750 230
rect 31990 -10 32080 230
rect 32320 -10 32410 230
rect 32650 -10 32740 230
rect 32980 -10 33070 230
rect 33310 -10 33400 230
rect 33640 -10 33730 230
rect 33970 -10 34060 230
rect 34300 -10 34390 230
rect 34630 -10 34720 230
rect 34960 -10 35050 230
rect 35290 -10 35460 230
rect 28520 -70 35460 -10
rect 28320 -100 35460 -70
rect 28320 -130 28780 -100
rect 28320 -200 28340 -130
rect 28410 -200 28450 -130
rect 28520 -200 28780 -130
rect 28320 -260 28780 -200
rect 28320 -330 28340 -260
rect 28410 -330 28450 -260
rect 28520 -330 28780 -260
rect 28320 -340 28780 -330
rect 29020 -340 29110 -100
rect 29350 -340 29440 -100
rect 29680 -340 29770 -100
rect 30010 -340 30100 -100
rect 30340 -340 30430 -100
rect 30670 -340 30760 -100
rect 31000 -340 31090 -100
rect 31330 -340 31420 -100
rect 31660 -340 31750 -100
rect 31990 -340 32080 -100
rect 32320 -340 32410 -100
rect 32650 -340 32740 -100
rect 32980 -340 33070 -100
rect 33310 -340 33400 -100
rect 33640 -340 33730 -100
rect 33970 -340 34060 -100
rect 34300 -340 34390 -100
rect 34630 -340 34720 -100
rect 34960 -340 35050 -100
rect 35290 -340 35460 -100
rect 28320 -350 35460 -340
rect 22320 -3160 28077 -3125
rect 22320 -3230 22340 -3160
rect 22410 -3230 22450 -3160
rect 22520 -3230 22560 -3160
rect 22630 -3230 28077 -3160
rect 22320 -3258 28077 -3230
rect 22320 -3270 22650 -3258
rect 22320 -3340 22340 -3270
rect 22410 -3340 22450 -3270
rect 22520 -3340 22560 -3270
rect 22630 -3340 22650 -3270
rect 22320 -3360 22650 -3340
rect 20020 -3690 20500 -3660
rect 20020 -3760 20070 -3690
rect 20470 -3760 20500 -3690
rect 20020 -3800 20080 -3760
rect 20450 -3800 20500 -3760
rect 20020 -3870 20070 -3800
rect 20470 -3870 20500 -3800
rect 20020 -3930 20080 -3870
rect 20450 -3930 20500 -3870
rect 20020 -3950 20500 -3930
rect 24500 -3690 24980 -3660
rect 24500 -3760 24550 -3690
rect 24950 -3760 24980 -3690
rect 24500 -3800 24560 -3760
rect 24930 -3800 24980 -3760
rect 24500 -3870 24550 -3800
rect 24950 -3870 24980 -3800
rect 24500 -3930 24560 -3870
rect 24930 -3930 24980 -3870
rect 24500 -3950 24980 -3930
rect 24000 -5890 24480 -5780
rect 24000 -5915 24110 -5890
rect 16575 -6025 24110 -5915
rect -2220 -6150 8490 -6130
rect -2220 -6220 8200 -6150
rect 8270 -6220 8300 -6150
rect 8370 -6220 8400 -6150
rect 8470 -6220 8490 -6150
rect -2220 -6250 8490 -6220
rect -2220 -6320 8200 -6250
rect 8270 -6320 8300 -6250
rect 8370 -6320 8400 -6250
rect 8470 -6320 8490 -6250
rect -2220 -6350 8490 -6320
rect -2220 -7870 -1940 -6350
rect -2220 -7940 -2200 -7870
rect -2130 -7940 -2090 -7870
rect -2020 -7940 -1940 -7870
rect -2220 -7980 -1940 -7940
rect -2220 -8050 -2200 -7980
rect -2130 -8050 -2090 -7980
rect -2020 -8050 -1940 -7980
rect -2220 -8090 -1940 -8050
rect -2220 -8160 -2200 -8090
rect -2130 -8160 -2090 -8090
rect -2020 -8160 -1940 -8090
rect -2220 -8200 -1940 -8160
rect -2220 -8270 -2200 -8200
rect -2130 -8270 -2090 -8200
rect -2020 -8270 -1940 -8200
rect -2220 -8290 -1940 -8270
rect -1860 -7660 -250 -7450
rect -1860 -7900 -1650 -7660
rect -1410 -7900 -1320 -7660
rect -1080 -7900 -990 -7660
rect -750 -7900 -660 -7660
rect -420 -7900 -250 -7660
rect -1860 -7990 -250 -7900
rect -1860 -8230 -1650 -7990
rect -1410 -8230 -1320 -7990
rect -1080 -8230 -990 -7990
rect -750 -8230 -660 -7990
rect -420 -8230 -250 -7990
rect -1860 -8320 -250 -8230
rect -1860 -8560 -1650 -8320
rect -1410 -8560 -1320 -8320
rect -1080 -8560 -990 -8320
rect -750 -8560 -660 -8320
rect -420 -8560 -250 -8320
rect -1860 -8580 -250 -8560
rect -2220 -8640 -250 -8580
rect -2220 -8710 -2140 -8640
rect -2070 -8710 -2030 -8640
rect -1960 -8650 -250 -8640
rect -1960 -8710 -1650 -8650
rect -2220 -8750 -1650 -8710
rect -2220 -8820 -2140 -8750
rect -2070 -8820 -2030 -8750
rect -1960 -8820 -1650 -8750
rect -2220 -8860 -1650 -8820
rect -2220 -8930 -2140 -8860
rect -2070 -8930 -2030 -8860
rect -1960 -8890 -1650 -8860
rect -1410 -8890 -1320 -8650
rect -1080 -8890 -990 -8650
rect -750 -8890 -660 -8650
rect -420 -8890 -250 -8650
rect -1960 -8930 -250 -8890
rect -170 -7630 150 -7620
rect -170 -7700 -160 -7630
rect -90 -7650 -70 -7630
rect 0 -7650 20 -7630
rect 90 -7650 150 -7630
rect -170 -7720 -120 -7700
rect -170 -7790 -160 -7720
rect -170 -7810 -120 -7790
rect -170 -7880 -160 -7810
rect -170 -7890 -120 -7880
rect 120 -7890 150 -7650
rect -170 -7900 150 -7890
rect -170 -7970 -160 -7900
rect -90 -7970 -70 -7900
rect 0 -7970 20 -7900
rect 90 -7970 150 -7900
rect -170 -7980 150 -7970
rect -170 -7990 -120 -7980
rect -170 -8060 -160 -7990
rect -170 -8080 -120 -8060
rect -170 -8150 -160 -8080
rect -170 -8170 -120 -8150
rect -170 -8240 -160 -8170
rect 120 -8220 150 -7980
rect -90 -8240 -70 -8220
rect 0 -8240 20 -8220
rect 90 -8230 150 -8220
rect 14590 -8230 14900 -8210
rect 90 -8240 9020 -8230
rect -170 -8250 9020 -8240
rect -170 -8260 8730 -8250
rect -170 -8330 -160 -8260
rect -90 -8310 -70 -8260
rect 0 -8310 20 -8260
rect 90 -8310 8730 -8260
rect 120 -8320 8730 -8310
rect 8800 -8320 8830 -8250
rect 8900 -8320 8930 -8250
rect 9000 -8320 9020 -8250
rect -170 -8350 -120 -8330
rect 120 -8350 9020 -8320
rect -170 -8420 -160 -8350
rect 120 -8420 8730 -8350
rect 8800 -8420 8830 -8350
rect 8900 -8420 8930 -8350
rect 9000 -8420 9020 -8350
rect -170 -8440 -120 -8420
rect 120 -8440 9020 -8420
rect 14590 -8300 14600 -8230
rect 14670 -8300 14700 -8230
rect 14770 -8300 14810 -8230
rect 14880 -8300 14900 -8230
rect 14590 -8325 14900 -8300
rect 16575 -8325 16685 -6025
rect 14590 -8340 16685 -8325
rect 14590 -8410 14600 -8340
rect 14670 -8410 14700 -8340
rect 14770 -8410 14810 -8340
rect 14880 -8410 16685 -8340
rect 14590 -8435 16685 -8410
rect -170 -8510 -160 -8440
rect -170 -8530 -120 -8510
rect -170 -8600 -160 -8530
rect 120 -8550 150 -8440
rect 14590 -8450 14900 -8435
rect 14590 -8520 14600 -8450
rect 14670 -8520 14700 -8450
rect 14770 -8520 14810 -8450
rect 14880 -8520 14900 -8450
rect 14590 -8540 14900 -8520
rect -90 -8600 -70 -8550
rect 0 -8600 20 -8550
rect 90 -8600 150 -8550
rect -170 -8620 150 -8600
rect -170 -8690 -160 -8620
rect -90 -8640 -70 -8620
rect 0 -8640 20 -8620
rect 90 -8640 150 -8620
rect -170 -8710 -120 -8690
rect -170 -8780 -160 -8710
rect -170 -8800 -120 -8780
rect -170 -8870 -160 -8800
rect -170 -8880 -120 -8870
rect 120 -8880 150 -8640
rect 19210 -8560 19530 -8530
rect 19210 -8630 19230 -8560
rect 19300 -8570 19330 -8560
rect 19400 -8570 19430 -8560
rect 19500 -8630 19530 -8560
rect 19210 -8660 19250 -8630
rect 19490 -8660 19530 -8630
rect 19210 -8730 19230 -8660
rect 19500 -8730 19530 -8660
rect 19210 -8760 19250 -8730
rect 19490 -8760 19530 -8730
rect 19210 -8830 19230 -8760
rect 19300 -8830 19330 -8810
rect 19400 -8830 19430 -8810
rect 19500 -8830 19530 -8760
rect 19210 -8850 19530 -8830
rect -170 -8910 150 -8880
rect -2220 -8970 -250 -8930
rect -2220 -9040 -2140 -8970
rect -2070 -9040 -2030 -8970
rect -1960 -9040 -250 -8970
rect -2220 -9060 -250 -9040
rect 19940 -9000 20260 -8970
rect 19940 -9070 19960 -9000
rect 20030 -9070 20060 -9000
rect 20130 -9070 20160 -9000
rect 20230 -9070 20260 -9000
rect 19940 -9100 20260 -9070
rect 19940 -9170 19960 -9100
rect 20030 -9170 20060 -9100
rect 20130 -9170 20160 -9100
rect 20230 -9170 20260 -9100
rect 19940 -9200 20260 -9170
rect 19940 -9270 19960 -9200
rect 20030 -9270 20060 -9200
rect 20130 -9270 20160 -9200
rect 20230 -9270 20260 -9200
rect 19940 -9390 20260 -9270
rect 1080 -10340 2680 -10310
rect 1080 -10410 1150 -10340
rect 1220 -10410 1260 -10340
rect 1550 -10410 1590 -10340
rect 1880 -10410 1920 -10340
rect 2210 -10410 2250 -10340
rect 2540 -10410 2580 -10340
rect 2650 -10410 2680 -10340
rect 1080 -10450 1260 -10410
rect 1500 -10450 1590 -10410
rect 1830 -10450 1930 -10410
rect 2170 -10450 2260 -10410
rect 2500 -10450 2680 -10410
rect 1080 -10520 1150 -10450
rect 1220 -10520 1260 -10450
rect 1550 -10520 1590 -10450
rect 1880 -10520 1920 -10450
rect 2210 -10520 2250 -10450
rect 2540 -10520 2580 -10450
rect 2650 -10520 2680 -10450
rect 1080 -10580 1260 -10520
rect 1500 -10580 1590 -10520
rect 1830 -10580 1930 -10520
rect 2170 -10580 2260 -10520
rect 2500 -10580 2680 -10520
rect 1080 -10600 2680 -10580
rect 12220 -10370 13820 -10340
rect 12220 -10440 12290 -10370
rect 12360 -10440 12400 -10370
rect 12690 -10440 12730 -10370
rect 13020 -10440 13060 -10370
rect 13350 -10440 13390 -10370
rect 13680 -10440 13720 -10370
rect 13790 -10440 13820 -10370
rect 12220 -10480 12400 -10440
rect 12640 -10480 12730 -10440
rect 12970 -10480 13070 -10440
rect 13310 -10480 13400 -10440
rect 13640 -10480 13820 -10440
rect 12220 -10550 12290 -10480
rect 12360 -10550 12400 -10480
rect 12690 -10550 12730 -10480
rect 13020 -10550 13060 -10480
rect 13350 -10550 13390 -10480
rect 13680 -10550 13720 -10480
rect 13790 -10550 13820 -10480
rect 12220 -10610 12400 -10550
rect 12640 -10610 12730 -10550
rect 12970 -10610 13070 -10550
rect 13310 -10610 13400 -10550
rect 13640 -10610 13820 -10550
rect 12220 -10620 13820 -10610
rect 27944 -10995 28077 -3258
rect 28700 -430 35460 -350
rect 28700 -670 28780 -430
rect 29020 -670 29110 -430
rect 29350 -670 29440 -430
rect 29680 -670 29770 -430
rect 30010 -670 30100 -430
rect 30340 -670 30430 -430
rect 30670 -670 30760 -430
rect 31000 -670 31090 -430
rect 31330 -670 31420 -430
rect 31660 -670 31750 -430
rect 31990 -670 32080 -430
rect 32320 -670 32410 -430
rect 32650 -670 32740 -430
rect 32980 -670 33070 -430
rect 33310 -670 33400 -430
rect 33640 -670 33730 -430
rect 33970 -670 34060 -430
rect 34300 -670 34390 -430
rect 34630 -670 34720 -430
rect 34960 -670 35050 -430
rect 35290 -670 35460 -430
rect 28700 -760 35460 -670
rect 28700 -1000 28780 -760
rect 29020 -1000 29110 -760
rect 29350 -1000 29440 -760
rect 29680 -1000 29770 -760
rect 30010 -1000 30100 -760
rect 30340 -1000 30430 -760
rect 30670 -1000 30760 -760
rect 31000 -1000 31090 -760
rect 31330 -1000 31420 -760
rect 31660 -1000 31750 -760
rect 31990 -1000 32080 -760
rect 32320 -1000 32410 -760
rect 32650 -1000 32740 -760
rect 32980 -1000 33070 -760
rect 33310 -1000 33400 -760
rect 33640 -1000 33730 -760
rect 33970 -1000 34060 -760
rect 34300 -1000 34390 -760
rect 34630 -1000 34720 -760
rect 34960 -1000 35050 -760
rect 35290 -1000 35460 -760
rect 28700 -1090 35460 -1000
rect 28700 -1330 28780 -1090
rect 29020 -1330 29110 -1090
rect 29350 -1330 29440 -1090
rect 29680 -1330 29770 -1090
rect 30010 -1330 30100 -1090
rect 30340 -1330 30430 -1090
rect 30670 -1330 30760 -1090
rect 31000 -1330 31090 -1090
rect 31330 -1330 31420 -1090
rect 31660 -1330 31750 -1090
rect 31990 -1330 32080 -1090
rect 32320 -1330 32410 -1090
rect 32650 -1330 32740 -1090
rect 32980 -1330 33070 -1090
rect 33310 -1330 33400 -1090
rect 33640 -1330 33730 -1090
rect 33970 -1330 34060 -1090
rect 34300 -1330 34390 -1090
rect 34630 -1330 34720 -1090
rect 34960 -1330 35050 -1090
rect 35290 -1330 35460 -1090
rect 28700 -1420 35460 -1330
rect 28700 -1660 28780 -1420
rect 29020 -1660 29110 -1420
rect 29350 -1660 29440 -1420
rect 29680 -1660 29770 -1420
rect 30010 -1660 30100 -1420
rect 30340 -1660 30430 -1420
rect 30670 -1660 30760 -1420
rect 31000 -1660 31090 -1420
rect 31330 -1660 31420 -1420
rect 31660 -1660 31750 -1420
rect 31990 -1660 32080 -1420
rect 32320 -1660 32410 -1420
rect 32650 -1660 32740 -1420
rect 32980 -1660 33070 -1420
rect 33310 -1660 33400 -1420
rect 33640 -1660 33730 -1420
rect 33970 -1660 34060 -1420
rect 34300 -1660 34390 -1420
rect 34630 -1660 34720 -1420
rect 34960 -1660 35050 -1420
rect 35290 -1660 35460 -1420
rect 28700 -1750 35460 -1660
rect 28700 -1990 28780 -1750
rect 29020 -1990 29110 -1750
rect 29350 -1990 29440 -1750
rect 29680 -1990 29770 -1750
rect 30010 -1990 30100 -1750
rect 30340 -1990 30430 -1750
rect 30670 -1990 30760 -1750
rect 31000 -1990 31090 -1750
rect 31330 -1990 31420 -1750
rect 31660 -1990 31750 -1750
rect 31990 -1990 32080 -1750
rect 32320 -1990 32410 -1750
rect 32650 -1990 32740 -1750
rect 32980 -1990 33070 -1750
rect 33310 -1990 33400 -1750
rect 33640 -1990 33730 -1750
rect 33970 -1990 34060 -1750
rect 34300 -1990 34390 -1750
rect 34630 -1990 34720 -1750
rect 34960 -1990 35050 -1750
rect 35290 -1990 35460 -1750
rect 28700 -2080 35460 -1990
rect 28700 -2320 28780 -2080
rect 29020 -2320 29110 -2080
rect 29350 -2320 29440 -2080
rect 29680 -2320 29770 -2080
rect 30010 -2320 30100 -2080
rect 30340 -2320 30430 -2080
rect 30670 -2320 30760 -2080
rect 31000 -2320 31090 -2080
rect 31330 -2320 31420 -2080
rect 31660 -2320 31750 -2080
rect 31990 -2320 32080 -2080
rect 32320 -2320 32410 -2080
rect 32650 -2320 32740 -2080
rect 32980 -2320 33070 -2080
rect 33310 -2320 33400 -2080
rect 33640 -2320 33730 -2080
rect 33970 -2320 34060 -2080
rect 34300 -2320 34390 -2080
rect 34630 -2320 34720 -2080
rect 34960 -2320 35050 -2080
rect 35290 -2320 35460 -2080
rect 28700 -2410 35460 -2320
rect 28700 -2650 28780 -2410
rect 29020 -2650 29110 -2410
rect 29350 -2650 29440 -2410
rect 29680 -2650 29770 -2410
rect 30010 -2650 30100 -2410
rect 30340 -2650 30430 -2410
rect 30670 -2650 30760 -2410
rect 31000 -2650 31090 -2410
rect 31330 -2650 31420 -2410
rect 31660 -2650 31750 -2410
rect 31990 -2650 32080 -2410
rect 32320 -2650 32410 -2410
rect 32650 -2650 32740 -2410
rect 32980 -2650 33070 -2410
rect 33310 -2650 33400 -2410
rect 33640 -2650 33730 -2410
rect 33970 -2650 34060 -2410
rect 34300 -2650 34390 -2410
rect 34630 -2650 34720 -2410
rect 34960 -2650 35050 -2410
rect 35290 -2650 35460 -2410
rect 28700 -2740 35460 -2650
rect 28700 -2980 28780 -2740
rect 29020 -2980 29110 -2740
rect 29350 -2980 29440 -2740
rect 29680 -2980 29770 -2740
rect 30010 -2980 30100 -2740
rect 30340 -2980 30430 -2740
rect 30670 -2980 30760 -2740
rect 31000 -2980 31090 -2740
rect 31330 -2980 31420 -2740
rect 31660 -2980 31750 -2740
rect 31990 -2980 32080 -2740
rect 32320 -2980 32410 -2740
rect 32650 -2980 32740 -2740
rect 32980 -2980 33070 -2740
rect 33310 -2980 33400 -2740
rect 33640 -2980 33730 -2740
rect 33970 -2980 34060 -2740
rect 34300 -2980 34390 -2740
rect 34630 -2980 34720 -2740
rect 34960 -2980 35050 -2740
rect 35290 -2980 35460 -2740
rect 28700 -3070 35460 -2980
rect 28700 -3310 28780 -3070
rect 29020 -3310 29110 -3070
rect 29350 -3310 29440 -3070
rect 29680 -3310 29770 -3070
rect 30010 -3310 30100 -3070
rect 30340 -3310 30430 -3070
rect 30670 -3310 30760 -3070
rect 31000 -3310 31090 -3070
rect 31330 -3310 31420 -3070
rect 31660 -3310 31750 -3070
rect 31990 -3310 32080 -3070
rect 32320 -3310 32410 -3070
rect 32650 -3310 32740 -3070
rect 32980 -3310 33070 -3070
rect 33310 -3310 33400 -3070
rect 33640 -3310 33730 -3070
rect 33970 -3310 34060 -3070
rect 34300 -3310 34390 -3070
rect 34630 -3310 34720 -3070
rect 34960 -3310 35050 -3070
rect 35290 -3310 35460 -3070
rect 28700 -3400 35460 -3310
rect 28700 -3640 28780 -3400
rect 29020 -3640 29110 -3400
rect 29350 -3640 29440 -3400
rect 29680 -3640 29770 -3400
rect 30010 -3640 30100 -3400
rect 30340 -3640 30430 -3400
rect 30670 -3640 30760 -3400
rect 31000 -3640 31090 -3400
rect 31330 -3640 31420 -3400
rect 31660 -3640 31750 -3400
rect 31990 -3640 32080 -3400
rect 32320 -3640 32410 -3400
rect 32650 -3640 32740 -3400
rect 32980 -3640 33070 -3400
rect 33310 -3640 33400 -3400
rect 33640 -3640 33730 -3400
rect 33970 -3640 34060 -3400
rect 34300 -3640 34390 -3400
rect 34630 -3640 34720 -3400
rect 34960 -3640 35050 -3400
rect 35290 -3640 35460 -3400
rect 28700 -3730 35460 -3640
rect 28700 -3970 28780 -3730
rect 29020 -3970 29110 -3730
rect 29350 -3970 29440 -3730
rect 29680 -3970 29770 -3730
rect 30010 -3970 30100 -3730
rect 30340 -3970 30430 -3730
rect 30670 -3970 30760 -3730
rect 31000 -3970 31090 -3730
rect 31330 -3970 31420 -3730
rect 31660 -3970 31750 -3730
rect 31990 -3970 32080 -3730
rect 32320 -3970 32410 -3730
rect 32650 -3970 32740 -3730
rect 32980 -3970 33070 -3730
rect 33310 -3970 33400 -3730
rect 33640 -3970 33730 -3730
rect 33970 -3970 34060 -3730
rect 34300 -3970 34390 -3730
rect 34630 -3970 34720 -3730
rect 34960 -3970 35050 -3730
rect 35290 -3970 35460 -3730
rect 28700 -4060 35460 -3970
rect 28700 -4300 28780 -4060
rect 29020 -4300 29110 -4060
rect 29350 -4300 29440 -4060
rect 29680 -4300 29770 -4060
rect 30010 -4300 30100 -4060
rect 30340 -4300 30430 -4060
rect 30670 -4300 30760 -4060
rect 31000 -4300 31090 -4060
rect 31330 -4300 31420 -4060
rect 31660 -4300 31750 -4060
rect 31990 -4300 32080 -4060
rect 32320 -4300 32410 -4060
rect 32650 -4300 32740 -4060
rect 32980 -4300 33070 -4060
rect 33310 -4300 33400 -4060
rect 33640 -4300 33730 -4060
rect 33970 -4300 34060 -4060
rect 34300 -4300 34390 -4060
rect 34630 -4300 34720 -4060
rect 34960 -4300 35050 -4060
rect 35290 -4300 35460 -4060
rect 28700 -4390 35460 -4300
rect 28700 -4630 28780 -4390
rect 29020 -4630 29110 -4390
rect 29350 -4630 29440 -4390
rect 29680 -4630 29770 -4390
rect 30010 -4630 30100 -4390
rect 30340 -4630 30430 -4390
rect 30670 -4630 30760 -4390
rect 31000 -4630 31090 -4390
rect 31330 -4630 31420 -4390
rect 31660 -4630 31750 -4390
rect 31990 -4630 32080 -4390
rect 32320 -4630 32410 -4390
rect 32650 -4630 32740 -4390
rect 32980 -4630 33070 -4390
rect 33310 -4630 33400 -4390
rect 33640 -4630 33730 -4390
rect 33970 -4630 34060 -4390
rect 34300 -4630 34390 -4390
rect 34630 -4630 34720 -4390
rect 34960 -4630 35050 -4390
rect 35290 -4630 35460 -4390
rect 28700 -4720 35460 -4630
rect 28700 -4960 28780 -4720
rect 29020 -4960 29110 -4720
rect 29350 -4960 29440 -4720
rect 29680 -4960 29770 -4720
rect 30010 -4960 30100 -4720
rect 30340 -4960 30430 -4720
rect 30670 -4960 30760 -4720
rect 31000 -4960 31090 -4720
rect 31330 -4960 31420 -4720
rect 31660 -4960 31750 -4720
rect 31990 -4960 32080 -4720
rect 32320 -4960 32410 -4720
rect 32650 -4960 32740 -4720
rect 32980 -4960 33070 -4720
rect 33310 -4960 33400 -4720
rect 33640 -4960 33730 -4720
rect 33970 -4960 34060 -4720
rect 34300 -4960 34390 -4720
rect 34630 -4960 34720 -4720
rect 34960 -4960 35050 -4720
rect 35290 -4960 35460 -4720
rect 28700 -5050 35460 -4960
rect 28700 -5290 28780 -5050
rect 29020 -5290 29110 -5050
rect 29350 -5290 29440 -5050
rect 29680 -5290 29770 -5050
rect 30010 -5290 30100 -5050
rect 30340 -5290 30430 -5050
rect 30670 -5290 30760 -5050
rect 31000 -5290 31090 -5050
rect 31330 -5290 31420 -5050
rect 31660 -5290 31750 -5050
rect 31990 -5290 32080 -5050
rect 32320 -5290 32410 -5050
rect 32650 -5290 32740 -5050
rect 32980 -5290 33070 -5050
rect 33310 -5290 33400 -5050
rect 33640 -5290 33730 -5050
rect 33970 -5290 34060 -5050
rect 34300 -5290 34390 -5050
rect 34630 -5290 34720 -5050
rect 34960 -5290 35050 -5050
rect 35290 -5290 35460 -5050
rect 28700 -5380 35460 -5290
rect 28700 -5620 28780 -5380
rect 29020 -5620 29110 -5380
rect 29350 -5620 29440 -5380
rect 29680 -5620 29770 -5380
rect 30010 -5620 30100 -5380
rect 30340 -5620 30430 -5380
rect 30670 -5620 30760 -5380
rect 31000 -5620 31090 -5380
rect 31330 -5620 31420 -5380
rect 31660 -5620 31750 -5380
rect 31990 -5620 32080 -5380
rect 32320 -5620 32410 -5380
rect 32650 -5620 32740 -5380
rect 32980 -5620 33070 -5380
rect 33310 -5620 33400 -5380
rect 33640 -5620 33730 -5380
rect 33970 -5620 34060 -5380
rect 34300 -5620 34390 -5380
rect 34630 -5620 34720 -5380
rect 34960 -5620 35050 -5380
rect 35290 -5620 35460 -5380
rect 28700 -5710 35460 -5620
rect 28700 -5950 28780 -5710
rect 29020 -5950 29110 -5710
rect 29350 -5950 29440 -5710
rect 29680 -5950 29770 -5710
rect 30010 -5950 30100 -5710
rect 30340 -5950 30430 -5710
rect 30670 -5950 30760 -5710
rect 31000 -5950 31090 -5710
rect 31330 -5950 31420 -5710
rect 31660 -5950 31750 -5710
rect 31990 -5950 32080 -5710
rect 32320 -5950 32410 -5710
rect 32650 -5950 32740 -5710
rect 32980 -5950 33070 -5710
rect 33310 -5950 33400 -5710
rect 33640 -5950 33730 -5710
rect 33970 -5950 34060 -5710
rect 34300 -5950 34390 -5710
rect 34630 -5950 34720 -5710
rect 34960 -5950 35050 -5710
rect 35290 -5950 35460 -5710
rect 28700 -6040 35460 -5950
rect 28700 -6280 28780 -6040
rect 29020 -6280 29110 -6040
rect 29350 -6280 29440 -6040
rect 29680 -6280 29770 -6040
rect 30010 -6280 30100 -6040
rect 30340 -6280 30430 -6040
rect 30670 -6280 30760 -6040
rect 31000 -6280 31090 -6040
rect 31330 -6280 31420 -6040
rect 31660 -6280 31750 -6040
rect 31990 -6280 32080 -6040
rect 32320 -6280 32410 -6040
rect 32650 -6280 32740 -6040
rect 32980 -6280 33070 -6040
rect 33310 -6280 33400 -6040
rect 33640 -6280 33730 -6040
rect 33970 -6280 34060 -6040
rect 34300 -6280 34390 -6040
rect 34630 -6280 34720 -6040
rect 34960 -6280 35050 -6040
rect 35290 -6280 35460 -6040
rect 28700 -6450 35460 -6280
rect 35780 220 36100 310
rect 35780 150 35790 220
rect 35860 170 35880 220
rect 35950 170 35970 220
rect 36040 170 36100 220
rect 35780 130 35830 150
rect 35780 60 35790 130
rect 35780 40 35830 60
rect 35780 -30 35790 40
rect 35780 -50 35830 -30
rect 35780 -120 35790 -50
rect 36070 -70 36100 170
rect 35860 -120 35880 -70
rect 35950 -120 35970 -70
rect 36040 -120 36100 -70
rect 35780 -140 36100 -120
rect 35780 -210 35790 -140
rect 35860 -160 35880 -140
rect 35950 -160 35970 -140
rect 36040 -160 36100 -140
rect 35780 -230 35830 -210
rect 35780 -300 35790 -230
rect 35780 -320 35830 -300
rect 35780 -390 35790 -320
rect 35780 -400 35830 -390
rect 36070 -400 36100 -160
rect 35780 -450 36100 -400
rect 35780 -520 35790 -450
rect 35860 -520 35880 -450
rect 35950 -520 35970 -450
rect 36040 -520 36100 -450
rect 35780 -530 36100 -520
rect 35780 -540 35830 -530
rect 35780 -610 35790 -540
rect 35780 -630 35830 -610
rect 35780 -700 35790 -630
rect 35780 -720 35830 -700
rect 35780 -790 35790 -720
rect 36070 -770 36100 -530
rect 35860 -790 35880 -770
rect 35950 -790 35970 -770
rect 36040 -790 36100 -770
rect 35780 -810 36100 -790
rect 35780 -880 35790 -810
rect 35860 -860 35880 -810
rect 35950 -860 35970 -810
rect 36040 -860 36100 -810
rect 35780 -900 35830 -880
rect 35780 -970 35790 -900
rect 35780 -990 35830 -970
rect 35780 -1060 35790 -990
rect 35780 -1080 35830 -1060
rect 35780 -1150 35790 -1080
rect 36070 -1100 36100 -860
rect 35860 -1150 35880 -1100
rect 35950 -1150 35970 -1100
rect 36040 -1150 36100 -1100
rect 35780 -1170 36100 -1150
rect 35780 -1240 35790 -1170
rect 35860 -1190 35880 -1170
rect 35950 -1190 35970 -1170
rect 36040 -1190 36100 -1170
rect 35780 -1260 35830 -1240
rect 35780 -1330 35790 -1260
rect 35780 -1350 35830 -1330
rect 35780 -1420 35790 -1350
rect 35780 -1430 35830 -1420
rect 36070 -1430 36100 -1190
rect 35780 -1440 36100 -1430
rect 35780 -1510 35790 -1440
rect 35860 -1510 35880 -1440
rect 35950 -1510 35970 -1440
rect 36040 -1510 36100 -1440
rect 35780 -1520 36100 -1510
rect 35780 -1530 35830 -1520
rect 35780 -1600 35790 -1530
rect 35780 -1620 35830 -1600
rect 35780 -1690 35790 -1620
rect 35780 -1710 35830 -1690
rect 35780 -1780 35790 -1710
rect 36070 -1760 36100 -1520
rect 35860 -1780 35880 -1760
rect 35950 -1780 35970 -1760
rect 36040 -1780 36100 -1760
rect 35780 -1800 36100 -1780
rect 35780 -1870 35790 -1800
rect 35860 -1850 35880 -1800
rect 35950 -1850 35970 -1800
rect 36040 -1850 36100 -1800
rect 35780 -1890 35830 -1870
rect 35780 -1960 35790 -1890
rect 35780 -1980 35830 -1960
rect 35780 -2050 35790 -1980
rect 35780 -2070 35830 -2050
rect 35780 -2140 35790 -2070
rect 36070 -2090 36100 -1850
rect 35860 -2140 35880 -2090
rect 35950 -2140 35970 -2090
rect 36040 -2140 36100 -2090
rect 35780 -2160 36100 -2140
rect 35780 -2230 35790 -2160
rect 35860 -2180 35880 -2160
rect 35950 -2180 35970 -2160
rect 36040 -2180 36100 -2160
rect 35780 -2250 35830 -2230
rect 35780 -2320 35790 -2250
rect 35780 -2340 35830 -2320
rect 35780 -2410 35790 -2340
rect 35780 -2420 35830 -2410
rect 36070 -2420 36100 -2180
rect 35780 -2430 36100 -2420
rect 35780 -2500 35790 -2430
rect 35860 -2500 35880 -2430
rect 35950 -2500 35970 -2430
rect 36040 -2500 36100 -2430
rect 35780 -2510 36100 -2500
rect 35780 -2520 35830 -2510
rect 35780 -2590 35790 -2520
rect 35780 -2610 35830 -2590
rect 35780 -2680 35790 -2610
rect 35780 -2700 35830 -2680
rect 35780 -2770 35790 -2700
rect 36070 -2750 36100 -2510
rect 35860 -2770 35880 -2750
rect 35950 -2770 35970 -2750
rect 36040 -2770 36100 -2750
rect 35780 -2790 36100 -2770
rect 35780 -2860 35790 -2790
rect 35860 -2840 35880 -2790
rect 35950 -2840 35970 -2790
rect 36040 -2840 36100 -2790
rect 35780 -2880 35830 -2860
rect 35780 -2950 35790 -2880
rect 35780 -2970 35830 -2950
rect 35780 -3040 35790 -2970
rect 35780 -3060 35830 -3040
rect 35780 -3130 35790 -3060
rect 36070 -3080 36100 -2840
rect 35860 -3130 35880 -3080
rect 35950 -3130 35970 -3080
rect 36040 -3130 36100 -3080
rect 35780 -3150 36100 -3130
rect 35780 -3220 35790 -3150
rect 35860 -3170 35880 -3150
rect 35950 -3170 35970 -3150
rect 36040 -3170 36100 -3150
rect 35780 -3240 35830 -3220
rect 35780 -3310 35790 -3240
rect 35780 -3330 35830 -3310
rect 35780 -3400 35790 -3330
rect 35780 -3410 35830 -3400
rect 36070 -3410 36100 -3170
rect 35780 -3460 36100 -3410
rect 35780 -3530 35790 -3460
rect 35860 -3530 35880 -3460
rect 35950 -3530 35970 -3460
rect 36040 -3530 36100 -3460
rect 35780 -3540 36100 -3530
rect 35780 -3550 35830 -3540
rect 35780 -3620 35790 -3550
rect 35780 -3640 35830 -3620
rect 35780 -3710 35790 -3640
rect 35780 -3730 35830 -3710
rect 35780 -3800 35790 -3730
rect 36070 -3780 36100 -3540
rect 35860 -3800 35880 -3780
rect 35950 -3800 35970 -3780
rect 36040 -3800 36100 -3780
rect 35780 -3820 36100 -3800
rect 35780 -3890 35790 -3820
rect 35860 -3870 35880 -3820
rect 35950 -3870 35970 -3820
rect 36040 -3870 36100 -3820
rect 35780 -3910 35830 -3890
rect 35780 -3980 35790 -3910
rect 35780 -4000 35830 -3980
rect 35780 -4070 35790 -4000
rect 35780 -4090 35830 -4070
rect 35780 -4160 35790 -4090
rect 36070 -4110 36100 -3870
rect 35860 -4160 35880 -4110
rect 35950 -4160 35970 -4110
rect 36040 -4160 36100 -4110
rect 35780 -4180 36100 -4160
rect 35780 -4250 35790 -4180
rect 35860 -4200 35880 -4180
rect 35950 -4200 35970 -4180
rect 36040 -4200 36100 -4180
rect 35780 -4270 35830 -4250
rect 35780 -4340 35790 -4270
rect 35780 -4360 35830 -4340
rect 35780 -4430 35790 -4360
rect 35780 -4440 35830 -4430
rect 36070 -4440 36100 -4200
rect 35780 -4450 36100 -4440
rect 35780 -4520 35790 -4450
rect 35860 -4520 35880 -4450
rect 35950 -4520 35970 -4450
rect 36040 -4520 36100 -4450
rect 35780 -4530 36100 -4520
rect 35780 -4540 35830 -4530
rect 35780 -4610 35790 -4540
rect 35780 -4630 35830 -4610
rect 35780 -4700 35790 -4630
rect 35780 -4720 35830 -4700
rect 35780 -4790 35790 -4720
rect 36070 -4770 36100 -4530
rect 35860 -4790 35880 -4770
rect 35950 -4790 35970 -4770
rect 36040 -4790 36100 -4770
rect 35780 -4810 36100 -4790
rect 35780 -4880 35790 -4810
rect 35860 -4860 35880 -4810
rect 35950 -4860 35970 -4810
rect 36040 -4860 36100 -4810
rect 35780 -4900 35830 -4880
rect 35780 -4970 35790 -4900
rect 35780 -4990 35830 -4970
rect 35780 -5060 35790 -4990
rect 35780 -5080 35830 -5060
rect 35780 -5150 35790 -5080
rect 36070 -5100 36100 -4860
rect 35860 -5150 35880 -5100
rect 35950 -5150 35970 -5100
rect 36040 -5150 36100 -5100
rect 35780 -5170 36100 -5150
rect 35780 -5240 35790 -5170
rect 35860 -5190 35880 -5170
rect 35950 -5190 35970 -5170
rect 36040 -5190 36100 -5170
rect 35780 -5260 35830 -5240
rect 35780 -5330 35790 -5260
rect 35780 -5350 35830 -5330
rect 35780 -5420 35790 -5350
rect 35780 -5430 35830 -5420
rect 36070 -5430 36100 -5190
rect 35780 -5440 36100 -5430
rect 35780 -5510 35790 -5440
rect 35860 -5510 35880 -5440
rect 35950 -5510 35970 -5440
rect 36040 -5510 36100 -5440
rect 35780 -5520 36100 -5510
rect 35780 -5530 35830 -5520
rect 35780 -5600 35790 -5530
rect 35780 -5620 35830 -5600
rect 35780 -5690 35790 -5620
rect 35780 -5710 35830 -5690
rect 35780 -5780 35790 -5710
rect 36070 -5760 36100 -5520
rect 35860 -5780 35880 -5760
rect 35950 -5780 35970 -5760
rect 36040 -5780 36100 -5760
rect 35780 -5800 36100 -5780
rect 35780 -5870 35790 -5800
rect 35860 -5850 35880 -5800
rect 35950 -5850 35970 -5800
rect 36040 -5850 36100 -5800
rect 35780 -5890 35830 -5870
rect 35780 -5960 35790 -5890
rect 35780 -5980 35830 -5960
rect 35780 -6050 35790 -5980
rect 35780 -6070 35830 -6050
rect 35780 -6140 35790 -6070
rect 36070 -6090 36100 -5850
rect 35860 -6140 35880 -6090
rect 35950 -6140 35970 -6090
rect 36040 -6140 36100 -6090
rect 35780 -6160 36100 -6140
rect 35780 -6230 35790 -6160
rect 35860 -6180 35880 -6160
rect 35950 -6180 35970 -6160
rect 36040 -6180 36100 -6160
rect 35780 -6250 35830 -6230
rect 35780 -6320 35790 -6250
rect 35780 -6340 35830 -6320
rect 35780 -6410 35790 -6340
rect 35780 -6420 35830 -6410
rect 36070 -6420 36100 -6180
rect 35780 -6450 36100 -6420
rect 24615 -11105 28077 -10995
rect 24615 -11600 24725 -11105
rect 24280 -11710 24760 -11600
rect 2210 -12240 3810 -12220
rect 2210 -12300 2390 -12240
rect 2630 -12300 2720 -12240
rect 2960 -12300 3060 -12240
rect 3300 -12300 3390 -12240
rect 3630 -12300 3810 -12240
rect 2210 -12370 2240 -12300
rect 2310 -12370 2350 -12300
rect 2640 -12370 2680 -12300
rect 2970 -12370 3010 -12300
rect 3300 -12370 3340 -12300
rect 3630 -12370 3670 -12300
rect 3740 -12370 3810 -12300
rect 2210 -12410 2390 -12370
rect 2630 -12410 2720 -12370
rect 2960 -12410 3060 -12370
rect 3300 -12410 3390 -12370
rect 3630 -12410 3810 -12370
rect 2210 -12480 2240 -12410
rect 2310 -12480 2350 -12410
rect 2640 -12480 2680 -12410
rect 2970 -12480 3010 -12410
rect 3300 -12480 3340 -12410
rect 3630 -12480 3670 -12410
rect 3740 -12480 3810 -12410
rect 2210 -12510 3810 -12480
rect 11090 -12240 12690 -12220
rect 11090 -12300 11270 -12240
rect 11510 -12300 11600 -12240
rect 11840 -12300 11940 -12240
rect 12180 -12300 12270 -12240
rect 12510 -12300 12690 -12240
rect 11090 -12370 11120 -12300
rect 11190 -12370 11230 -12300
rect 11520 -12370 11560 -12300
rect 11850 -12370 11890 -12300
rect 12180 -12370 12220 -12300
rect 12510 -12370 12550 -12300
rect 12620 -12370 12690 -12300
rect 11090 -12410 11270 -12370
rect 11510 -12410 11600 -12370
rect 11840 -12410 11940 -12370
rect 12180 -12410 12270 -12370
rect 12510 -12410 12690 -12370
rect 11090 -12480 11120 -12410
rect 11190 -12480 11230 -12410
rect 11520 -12480 11560 -12410
rect 11850 -12480 11890 -12410
rect 12180 -12480 12220 -12410
rect 12510 -12480 12550 -12410
rect 12620 -12480 12690 -12410
rect 11090 -12510 12690 -12480
rect 19210 -14220 19530 -14190
rect 19210 -14290 19230 -14220
rect 19300 -14230 19330 -14220
rect 19400 -14230 19430 -14220
rect 19500 -14290 19530 -14220
rect 19210 -14320 19250 -14290
rect 19490 -14320 19530 -14290
rect 19210 -14390 19230 -14320
rect 19500 -14390 19530 -14320
rect 19210 -14420 19250 -14390
rect 19490 -14420 19530 -14390
rect 19210 -14490 19230 -14420
rect 19300 -14490 19330 -14470
rect 19400 -14490 19430 -14470
rect 19500 -14490 19530 -14420
rect 19210 -14510 19530 -14490
rect 20460 -14870 20780 -14840
rect 20460 -14940 20480 -14870
rect 20550 -14940 20580 -14870
rect 20650 -14940 20680 -14870
rect 20750 -14940 20780 -14870
rect 20460 -14970 20780 -14940
rect 20460 -15040 20480 -14970
rect 20550 -15040 20580 -14970
rect 20650 -15040 20680 -14970
rect 20750 -15040 20780 -14970
rect 20460 -15070 20780 -15040
rect 20460 -15140 20480 -15070
rect 20550 -15140 20580 -15070
rect 20650 -15140 20680 -15070
rect 20750 -15140 20780 -15070
rect 20460 -15260 20780 -15140
rect 7210 -17600 7650 -17580
rect 7210 -17670 7230 -17600
rect 7300 -17670 7340 -17600
rect 7410 -17670 7450 -17600
rect 7520 -17670 7560 -17600
rect 7630 -17670 7650 -17600
rect 7210 -17680 7650 -17670
rect 24080 -17620 24560 -17500
rect 24080 -17680 24200 -17620
rect 7210 -17710 24200 -17680
rect 7210 -17780 7230 -17710
rect 7300 -17780 7340 -17710
rect 7410 -17780 7450 -17710
rect 7520 -17780 7560 -17710
rect 7630 -17780 24200 -17710
rect 7210 -17800 24200 -17780
rect 7210 -17820 7650 -17800
rect 7210 -17890 7230 -17820
rect 7300 -17890 7340 -17820
rect 7410 -17890 7450 -17820
rect 7520 -17890 7560 -17820
rect 7630 -17890 7650 -17820
rect 7210 -17930 7650 -17890
rect 7210 -18000 7230 -17930
rect 7300 -18000 7340 -17930
rect 7410 -18000 7450 -17930
rect 7520 -18000 7560 -17930
rect 7630 -18000 7650 -17930
rect 7210 -18020 7650 -18000
rect 19210 -20290 19530 -20260
rect 19210 -20360 19230 -20290
rect 19300 -20300 19330 -20290
rect 19400 -20300 19430 -20290
rect 19500 -20360 19530 -20290
rect 19210 -20390 19250 -20360
rect 19490 -20390 19530 -20360
rect 19210 -20460 19230 -20390
rect 19500 -20460 19530 -20390
rect 19210 -20490 19250 -20460
rect 19490 -20490 19530 -20460
rect 19210 -20560 19230 -20490
rect 19300 -20560 19330 -20540
rect 19400 -20560 19430 -20540
rect 19500 -20560 19530 -20490
rect 19210 -20580 19530 -20560
rect 20020 -20720 20340 -20690
rect 20020 -20790 20040 -20720
rect 20110 -20790 20140 -20720
rect 20210 -20790 20240 -20720
rect 20310 -20790 20340 -20720
rect 20020 -20820 20340 -20790
rect 20020 -20890 20040 -20820
rect 20110 -20890 20140 -20820
rect 20210 -20890 20240 -20820
rect 20310 -20890 20340 -20820
rect 20020 -20920 20340 -20890
rect 20020 -20990 20040 -20920
rect 20110 -20990 20140 -20920
rect 20210 -20990 20240 -20920
rect 20310 -20990 20340 -20920
rect 20020 -21110 20340 -20990
rect 2210 -22660 3810 -22630
rect 2210 -22730 2280 -22660
rect 2350 -22730 2390 -22660
rect 2680 -22730 2720 -22660
rect 3010 -22730 3050 -22660
rect 3340 -22730 3380 -22660
rect 3670 -22730 3710 -22660
rect 3780 -22730 3810 -22660
rect 2210 -22770 2390 -22730
rect 2630 -22770 2720 -22730
rect 2960 -22770 3060 -22730
rect 3300 -22770 3390 -22730
rect 3630 -22770 3810 -22730
rect 2210 -22840 2280 -22770
rect 2350 -22840 2390 -22770
rect 2680 -22840 2720 -22770
rect 3010 -22840 3050 -22770
rect 3340 -22840 3380 -22770
rect 3670 -22840 3710 -22770
rect 3780 -22840 3810 -22770
rect 2210 -22900 2390 -22840
rect 2630 -22900 2720 -22840
rect 2960 -22900 3060 -22840
rect 3300 -22900 3390 -22840
rect 3630 -22900 3810 -22840
rect 2210 -22910 3810 -22900
rect 11090 -22660 12690 -22630
rect 11090 -22730 11160 -22660
rect 11230 -22730 11270 -22660
rect 11560 -22730 11600 -22660
rect 11890 -22730 11930 -22660
rect 12220 -22730 12260 -22660
rect 12550 -22730 12590 -22660
rect 12660 -22730 12690 -22660
rect 11090 -22770 11270 -22730
rect 11510 -22770 11600 -22730
rect 11840 -22770 11940 -22730
rect 12180 -22770 12270 -22730
rect 12510 -22770 12690 -22730
rect 11090 -22840 11160 -22770
rect 11230 -22840 11270 -22770
rect 11560 -22840 11600 -22770
rect 11890 -22840 11930 -22770
rect 12220 -22840 12260 -22770
rect 12550 -22840 12590 -22770
rect 12660 -22840 12690 -22770
rect 11090 -22900 11270 -22840
rect 11510 -22900 11600 -22840
rect 11840 -22900 11940 -22840
rect 12180 -22900 12270 -22840
rect 12510 -22900 12690 -22840
rect 11090 -22910 12690 -22900
<< via4 >>
rect -4650 8430 -4640 8460
rect -4640 8430 -4570 8460
rect -4570 8430 -4550 8460
rect -4550 8430 -4480 8460
rect -4480 8430 -4460 8460
rect -4460 8430 -4410 8460
rect -4320 8430 -4300 8460
rect -4300 8430 -4280 8460
rect -4280 8430 -4210 8460
rect -4210 8430 -4190 8460
rect -4190 8430 -4120 8460
rect -4120 8430 -4100 8460
rect -4100 8430 -4080 8460
rect -3990 8430 -3940 8460
rect -3940 8430 -3920 8460
rect -3920 8430 -3850 8460
rect -3850 8430 -3830 8460
rect -3830 8430 -3760 8460
rect -3760 8430 -3750 8460
rect -3660 8430 -3650 8460
rect -3650 8430 -3580 8460
rect -3580 8430 -3560 8460
rect -3560 8430 -3490 8460
rect -3490 8430 -3470 8460
rect -3470 8430 -3420 8460
rect -3330 8430 -3310 8460
rect -3310 8430 -3290 8460
rect -3290 8430 -3220 8460
rect -3220 8430 -3200 8460
rect -3200 8430 -3130 8460
rect -3130 8430 -3110 8460
rect -3110 8430 -3090 8460
rect -3000 8430 -2950 8460
rect -2950 8430 -2930 8460
rect -2930 8430 -2860 8460
rect -2860 8430 -2840 8460
rect -2840 8430 -2770 8460
rect -2770 8430 -2760 8460
rect -2670 8430 -2660 8460
rect -2660 8430 -2590 8460
rect -2590 8430 -2570 8460
rect -2570 8430 -2500 8460
rect -2500 8430 -2480 8460
rect -2480 8430 -2430 8460
rect -2340 8430 -2320 8460
rect -2320 8430 -2300 8460
rect -2300 8430 -2230 8460
rect -2230 8430 -2210 8460
rect -2210 8430 -2140 8460
rect -2140 8430 -2120 8460
rect -2120 8430 -2100 8460
rect -2010 8430 -1960 8460
rect -1960 8430 -1940 8460
rect -1940 8430 -1870 8460
rect -1870 8430 -1850 8460
rect -1850 8430 -1780 8460
rect -1780 8430 -1770 8460
rect -1640 8430 -1630 8460
rect -1630 8430 -1560 8460
rect -1560 8430 -1540 8460
rect -1540 8430 -1470 8460
rect -1470 8430 -1450 8460
rect -1450 8430 -1400 8460
rect -1310 8430 -1290 8460
rect -1290 8430 -1270 8460
rect -1270 8430 -1200 8460
rect -1200 8430 -1180 8460
rect -1180 8430 -1110 8460
rect -1110 8430 -1090 8460
rect -1090 8430 -1070 8460
rect -980 8430 -930 8460
rect -930 8430 -910 8460
rect -910 8430 -840 8460
rect -840 8430 -820 8460
rect -820 8430 -750 8460
rect -750 8430 -740 8460
rect -650 8430 -640 8460
rect -640 8430 -570 8460
rect -570 8430 -550 8460
rect -550 8430 -480 8460
rect -480 8430 -460 8460
rect -460 8430 -410 8460
rect -320 8430 -300 8460
rect -300 8430 -280 8460
rect -280 8430 -210 8460
rect -210 8430 -190 8460
rect -190 8430 -120 8460
rect -120 8430 -100 8460
rect -100 8430 -80 8460
rect 10 8430 60 8460
rect 60 8430 80 8460
rect 80 8430 150 8460
rect 150 8430 170 8460
rect 170 8430 240 8460
rect 240 8430 250 8460
rect 340 8430 350 8460
rect 350 8430 420 8460
rect 420 8430 440 8460
rect 440 8430 510 8460
rect 510 8430 530 8460
rect 530 8430 580 8460
rect 670 8430 690 8460
rect 690 8430 710 8460
rect 710 8430 780 8460
rect 780 8430 800 8460
rect 800 8430 870 8460
rect 870 8430 890 8460
rect 890 8430 910 8460
rect 1000 8430 1050 8460
rect 1050 8430 1070 8460
rect 1070 8430 1140 8460
rect 1140 8430 1160 8460
rect 1160 8430 1230 8460
rect 1230 8430 1240 8460
rect 1370 8430 1380 8460
rect 1380 8430 1450 8460
rect 1450 8430 1470 8460
rect 1470 8430 1540 8460
rect 1540 8430 1560 8460
rect 1560 8430 1610 8460
rect 1700 8430 1720 8460
rect 1720 8430 1740 8460
rect 1740 8430 1810 8460
rect 1810 8430 1830 8460
rect 1830 8430 1900 8460
rect 1900 8430 1920 8460
rect 1920 8430 1940 8460
rect 2030 8430 2080 8460
rect 2080 8430 2100 8460
rect 2100 8430 2170 8460
rect 2170 8430 2190 8460
rect 2190 8430 2260 8460
rect 2260 8430 2270 8460
rect 2360 8430 2370 8460
rect 2370 8430 2440 8460
rect 2440 8430 2460 8460
rect 2460 8430 2530 8460
rect 2530 8430 2550 8460
rect 2550 8430 2600 8460
rect 2690 8430 2710 8460
rect 2710 8430 2730 8460
rect 2730 8430 2800 8460
rect 2800 8430 2820 8460
rect 2820 8430 2890 8460
rect 2890 8430 2910 8460
rect 2910 8430 2930 8460
rect 3020 8430 3070 8460
rect 3070 8430 3090 8460
rect 3090 8430 3160 8460
rect 3160 8430 3180 8460
rect 3180 8430 3250 8460
rect 3250 8430 3260 8460
rect 3350 8430 3360 8460
rect 3360 8430 3430 8460
rect 3430 8430 3450 8460
rect 3450 8430 3520 8460
rect 3520 8430 3540 8460
rect 3540 8430 3590 8460
rect 3680 8430 3700 8460
rect 3700 8430 3720 8460
rect 3720 8430 3790 8460
rect 3790 8430 3810 8460
rect 3810 8430 3880 8460
rect 3880 8430 3900 8460
rect 3900 8430 3920 8460
rect 4010 8430 4060 8460
rect 4060 8430 4080 8460
rect 4080 8430 4150 8460
rect 4150 8430 4170 8460
rect 4170 8430 4240 8460
rect 4240 8430 4250 8460
rect 4380 8430 4390 8460
rect 4390 8430 4460 8460
rect 4460 8430 4480 8460
rect 4480 8430 4550 8460
rect 4550 8430 4570 8460
rect 4570 8430 4620 8460
rect 4710 8430 4730 8460
rect 4730 8430 4750 8460
rect 4750 8430 4820 8460
rect 4820 8430 4840 8460
rect 4840 8430 4910 8460
rect 4910 8430 4930 8460
rect 4930 8430 4950 8460
rect 5040 8430 5090 8460
rect 5090 8430 5110 8460
rect 5110 8430 5180 8460
rect 5180 8430 5200 8460
rect 5200 8430 5270 8460
rect 5270 8430 5280 8460
rect 5370 8430 5380 8460
rect 5380 8430 5450 8460
rect 5450 8430 5470 8460
rect 5470 8430 5540 8460
rect 5540 8430 5560 8460
rect 5560 8430 5610 8460
rect 5700 8430 5720 8460
rect 5720 8430 5740 8460
rect 5740 8430 5810 8460
rect 5810 8430 5830 8460
rect 5830 8430 5900 8460
rect 5900 8430 5920 8460
rect 5920 8430 5940 8460
rect 6030 8430 6080 8460
rect 6080 8430 6100 8460
rect 6100 8430 6170 8460
rect 6170 8430 6190 8460
rect 6190 8430 6260 8460
rect 6260 8430 6270 8460
rect 6360 8430 6370 8460
rect 6370 8430 6440 8460
rect 6440 8430 6460 8460
rect 6460 8430 6530 8460
rect 6530 8430 6550 8460
rect 6550 8430 6600 8460
rect 6690 8430 6710 8460
rect 6710 8430 6730 8460
rect 6730 8430 6800 8460
rect 6800 8430 6820 8460
rect 6820 8430 6890 8460
rect 6890 8430 6910 8460
rect 6910 8430 6930 8460
rect 7020 8430 7070 8460
rect 7070 8430 7090 8460
rect 7090 8430 7160 8460
rect 7160 8430 7180 8460
rect 7180 8430 7250 8460
rect 7250 8430 7260 8460
rect -4650 8410 -4410 8430
rect -4320 8410 -4080 8430
rect -3990 8410 -3750 8430
rect -3660 8410 -3420 8430
rect -3330 8410 -3090 8430
rect -3000 8410 -2760 8430
rect -2670 8410 -2430 8430
rect -2340 8410 -2100 8430
rect -2010 8410 -1770 8430
rect -1640 8410 -1400 8430
rect -1310 8410 -1070 8430
rect -980 8410 -740 8430
rect -650 8410 -410 8430
rect -320 8410 -80 8430
rect 10 8410 250 8430
rect 340 8410 580 8430
rect 670 8410 910 8430
rect 1000 8410 1240 8430
rect 1370 8410 1610 8430
rect 1700 8410 1940 8430
rect 2030 8410 2270 8430
rect 2360 8410 2600 8430
rect 2690 8410 2930 8430
rect 3020 8410 3260 8430
rect 3350 8410 3590 8430
rect 3680 8410 3920 8430
rect 4010 8410 4250 8430
rect 4380 8410 4620 8430
rect 4710 8410 4950 8430
rect 5040 8410 5280 8430
rect 5370 8410 5610 8430
rect 5700 8410 5940 8430
rect 6030 8410 6270 8430
rect 6360 8410 6600 8430
rect 6690 8410 6930 8430
rect 7020 8410 7260 8430
rect -4650 8340 -4640 8410
rect -4640 8340 -4570 8410
rect -4570 8340 -4550 8410
rect -4550 8340 -4480 8410
rect -4480 8340 -4460 8410
rect -4460 8340 -4410 8410
rect -4320 8340 -4300 8410
rect -4300 8340 -4280 8410
rect -4280 8340 -4210 8410
rect -4210 8340 -4190 8410
rect -4190 8340 -4120 8410
rect -4120 8340 -4100 8410
rect -4100 8340 -4080 8410
rect -3990 8340 -3940 8410
rect -3940 8340 -3920 8410
rect -3920 8340 -3850 8410
rect -3850 8340 -3830 8410
rect -3830 8340 -3760 8410
rect -3760 8340 -3750 8410
rect -3660 8340 -3650 8410
rect -3650 8340 -3580 8410
rect -3580 8340 -3560 8410
rect -3560 8340 -3490 8410
rect -3490 8340 -3470 8410
rect -3470 8340 -3420 8410
rect -3330 8340 -3310 8410
rect -3310 8340 -3290 8410
rect -3290 8340 -3220 8410
rect -3220 8340 -3200 8410
rect -3200 8340 -3130 8410
rect -3130 8340 -3110 8410
rect -3110 8340 -3090 8410
rect -3000 8340 -2950 8410
rect -2950 8340 -2930 8410
rect -2930 8340 -2860 8410
rect -2860 8340 -2840 8410
rect -2840 8340 -2770 8410
rect -2770 8340 -2760 8410
rect -2670 8340 -2660 8410
rect -2660 8340 -2590 8410
rect -2590 8340 -2570 8410
rect -2570 8340 -2500 8410
rect -2500 8340 -2480 8410
rect -2480 8340 -2430 8410
rect -2340 8340 -2320 8410
rect -2320 8340 -2300 8410
rect -2300 8340 -2230 8410
rect -2230 8340 -2210 8410
rect -2210 8340 -2140 8410
rect -2140 8340 -2120 8410
rect -2120 8340 -2100 8410
rect -2010 8340 -1960 8410
rect -1960 8340 -1940 8410
rect -1940 8340 -1870 8410
rect -1870 8340 -1850 8410
rect -1850 8340 -1780 8410
rect -1780 8340 -1770 8410
rect -1640 8340 -1630 8410
rect -1630 8340 -1560 8410
rect -1560 8340 -1540 8410
rect -1540 8340 -1470 8410
rect -1470 8340 -1450 8410
rect -1450 8340 -1400 8410
rect -1310 8340 -1290 8410
rect -1290 8340 -1270 8410
rect -1270 8340 -1200 8410
rect -1200 8340 -1180 8410
rect -1180 8340 -1110 8410
rect -1110 8340 -1090 8410
rect -1090 8340 -1070 8410
rect -980 8340 -930 8410
rect -930 8340 -910 8410
rect -910 8340 -840 8410
rect -840 8340 -820 8410
rect -820 8340 -750 8410
rect -750 8340 -740 8410
rect -650 8340 -640 8410
rect -640 8340 -570 8410
rect -570 8340 -550 8410
rect -550 8340 -480 8410
rect -480 8340 -460 8410
rect -460 8340 -410 8410
rect -320 8340 -300 8410
rect -300 8340 -280 8410
rect -280 8340 -210 8410
rect -210 8340 -190 8410
rect -190 8340 -120 8410
rect -120 8340 -100 8410
rect -100 8340 -80 8410
rect 10 8340 60 8410
rect 60 8340 80 8410
rect 80 8340 150 8410
rect 150 8340 170 8410
rect 170 8340 240 8410
rect 240 8340 250 8410
rect 340 8340 350 8410
rect 350 8340 420 8410
rect 420 8340 440 8410
rect 440 8340 510 8410
rect 510 8340 530 8410
rect 530 8340 580 8410
rect 670 8340 690 8410
rect 690 8340 710 8410
rect 710 8340 780 8410
rect 780 8340 800 8410
rect 800 8340 870 8410
rect 870 8340 890 8410
rect 890 8340 910 8410
rect 1000 8340 1050 8410
rect 1050 8340 1070 8410
rect 1070 8340 1140 8410
rect 1140 8340 1160 8410
rect 1160 8340 1230 8410
rect 1230 8340 1240 8410
rect 1370 8340 1380 8410
rect 1380 8340 1450 8410
rect 1450 8340 1470 8410
rect 1470 8340 1540 8410
rect 1540 8340 1560 8410
rect 1560 8340 1610 8410
rect 1700 8340 1720 8410
rect 1720 8340 1740 8410
rect 1740 8340 1810 8410
rect 1810 8340 1830 8410
rect 1830 8340 1900 8410
rect 1900 8340 1920 8410
rect 1920 8340 1940 8410
rect 2030 8340 2080 8410
rect 2080 8340 2100 8410
rect 2100 8340 2170 8410
rect 2170 8340 2190 8410
rect 2190 8340 2260 8410
rect 2260 8340 2270 8410
rect 2360 8340 2370 8410
rect 2370 8340 2440 8410
rect 2440 8340 2460 8410
rect 2460 8340 2530 8410
rect 2530 8340 2550 8410
rect 2550 8340 2600 8410
rect 2690 8340 2710 8410
rect 2710 8340 2730 8410
rect 2730 8340 2800 8410
rect 2800 8340 2820 8410
rect 2820 8340 2890 8410
rect 2890 8340 2910 8410
rect 2910 8340 2930 8410
rect 3020 8340 3070 8410
rect 3070 8340 3090 8410
rect 3090 8340 3160 8410
rect 3160 8340 3180 8410
rect 3180 8340 3250 8410
rect 3250 8340 3260 8410
rect 3350 8340 3360 8410
rect 3360 8340 3430 8410
rect 3430 8340 3450 8410
rect 3450 8340 3520 8410
rect 3520 8340 3540 8410
rect 3540 8340 3590 8410
rect 3680 8340 3700 8410
rect 3700 8340 3720 8410
rect 3720 8340 3790 8410
rect 3790 8340 3810 8410
rect 3810 8340 3880 8410
rect 3880 8340 3900 8410
rect 3900 8340 3920 8410
rect 4010 8340 4060 8410
rect 4060 8340 4080 8410
rect 4080 8340 4150 8410
rect 4150 8340 4170 8410
rect 4170 8340 4240 8410
rect 4240 8340 4250 8410
rect 4380 8340 4390 8410
rect 4390 8340 4460 8410
rect 4460 8340 4480 8410
rect 4480 8340 4550 8410
rect 4550 8340 4570 8410
rect 4570 8340 4620 8410
rect 4710 8340 4730 8410
rect 4730 8340 4750 8410
rect 4750 8340 4820 8410
rect 4820 8340 4840 8410
rect 4840 8340 4910 8410
rect 4910 8340 4930 8410
rect 4930 8340 4950 8410
rect 5040 8340 5090 8410
rect 5090 8340 5110 8410
rect 5110 8340 5180 8410
rect 5180 8340 5200 8410
rect 5200 8340 5270 8410
rect 5270 8340 5280 8410
rect 5370 8340 5380 8410
rect 5380 8340 5450 8410
rect 5450 8340 5470 8410
rect 5470 8340 5540 8410
rect 5540 8340 5560 8410
rect 5560 8340 5610 8410
rect 5700 8340 5720 8410
rect 5720 8340 5740 8410
rect 5740 8340 5810 8410
rect 5810 8340 5830 8410
rect 5830 8340 5900 8410
rect 5900 8340 5920 8410
rect 5920 8340 5940 8410
rect 6030 8340 6080 8410
rect 6080 8340 6100 8410
rect 6100 8340 6170 8410
rect 6170 8340 6190 8410
rect 6190 8340 6260 8410
rect 6260 8340 6270 8410
rect 6360 8340 6370 8410
rect 6370 8340 6440 8410
rect 6440 8340 6460 8410
rect 6460 8340 6530 8410
rect 6530 8340 6550 8410
rect 6550 8340 6600 8410
rect 6690 8340 6710 8410
rect 6710 8340 6730 8410
rect 6730 8340 6800 8410
rect 6800 8340 6820 8410
rect 6820 8340 6890 8410
rect 6890 8340 6910 8410
rect 6910 8340 6930 8410
rect 7020 8340 7070 8410
rect 7070 8340 7090 8410
rect 7090 8340 7160 8410
rect 7160 8340 7180 8410
rect 7180 8340 7250 8410
rect 7250 8340 7260 8410
rect -4650 8320 -4410 8340
rect -4320 8320 -4080 8340
rect -3990 8320 -3750 8340
rect -3660 8320 -3420 8340
rect -3330 8320 -3090 8340
rect -3000 8320 -2760 8340
rect -2670 8320 -2430 8340
rect -2340 8320 -2100 8340
rect -2010 8320 -1770 8340
rect -1640 8320 -1400 8340
rect -1310 8320 -1070 8340
rect -980 8320 -740 8340
rect -650 8320 -410 8340
rect -320 8320 -80 8340
rect 10 8320 250 8340
rect 340 8320 580 8340
rect 670 8320 910 8340
rect 1000 8320 1240 8340
rect 1370 8320 1610 8340
rect 1700 8320 1940 8340
rect 2030 8320 2270 8340
rect 2360 8320 2600 8340
rect 2690 8320 2930 8340
rect 3020 8320 3260 8340
rect 3350 8320 3590 8340
rect 3680 8320 3920 8340
rect 4010 8320 4250 8340
rect 4380 8320 4620 8340
rect 4710 8320 4950 8340
rect 5040 8320 5280 8340
rect 5370 8320 5610 8340
rect 5700 8320 5940 8340
rect 6030 8320 6270 8340
rect 6360 8320 6600 8340
rect 6690 8320 6930 8340
rect 7020 8320 7260 8340
rect -4650 8250 -4640 8320
rect -4640 8250 -4570 8320
rect -4570 8250 -4550 8320
rect -4550 8250 -4480 8320
rect -4480 8250 -4460 8320
rect -4460 8250 -4410 8320
rect -4320 8250 -4300 8320
rect -4300 8250 -4280 8320
rect -4280 8250 -4210 8320
rect -4210 8250 -4190 8320
rect -4190 8250 -4120 8320
rect -4120 8250 -4100 8320
rect -4100 8250 -4080 8320
rect -3990 8250 -3940 8320
rect -3940 8250 -3920 8320
rect -3920 8250 -3850 8320
rect -3850 8250 -3830 8320
rect -3830 8250 -3760 8320
rect -3760 8250 -3750 8320
rect -3660 8250 -3650 8320
rect -3650 8250 -3580 8320
rect -3580 8250 -3560 8320
rect -3560 8250 -3490 8320
rect -3490 8250 -3470 8320
rect -3470 8250 -3420 8320
rect -3330 8250 -3310 8320
rect -3310 8250 -3290 8320
rect -3290 8250 -3220 8320
rect -3220 8250 -3200 8320
rect -3200 8250 -3130 8320
rect -3130 8250 -3110 8320
rect -3110 8250 -3090 8320
rect -3000 8250 -2950 8320
rect -2950 8250 -2930 8320
rect -2930 8250 -2860 8320
rect -2860 8250 -2840 8320
rect -2840 8250 -2770 8320
rect -2770 8250 -2760 8320
rect -2670 8250 -2660 8320
rect -2660 8250 -2590 8320
rect -2590 8250 -2570 8320
rect -2570 8250 -2500 8320
rect -2500 8250 -2480 8320
rect -2480 8250 -2430 8320
rect -2340 8250 -2320 8320
rect -2320 8250 -2300 8320
rect -2300 8250 -2230 8320
rect -2230 8250 -2210 8320
rect -2210 8250 -2140 8320
rect -2140 8250 -2120 8320
rect -2120 8250 -2100 8320
rect -2010 8250 -1960 8320
rect -1960 8250 -1940 8320
rect -1940 8250 -1870 8320
rect -1870 8250 -1850 8320
rect -1850 8250 -1780 8320
rect -1780 8250 -1770 8320
rect -1640 8250 -1630 8320
rect -1630 8250 -1560 8320
rect -1560 8250 -1540 8320
rect -1540 8250 -1470 8320
rect -1470 8250 -1450 8320
rect -1450 8250 -1400 8320
rect -1310 8250 -1290 8320
rect -1290 8250 -1270 8320
rect -1270 8250 -1200 8320
rect -1200 8250 -1180 8320
rect -1180 8250 -1110 8320
rect -1110 8250 -1090 8320
rect -1090 8250 -1070 8320
rect -980 8250 -930 8320
rect -930 8250 -910 8320
rect -910 8250 -840 8320
rect -840 8250 -820 8320
rect -820 8250 -750 8320
rect -750 8250 -740 8320
rect -650 8250 -640 8320
rect -640 8250 -570 8320
rect -570 8250 -550 8320
rect -550 8250 -480 8320
rect -480 8250 -460 8320
rect -460 8250 -410 8320
rect -320 8250 -300 8320
rect -300 8250 -280 8320
rect -280 8250 -210 8320
rect -210 8250 -190 8320
rect -190 8250 -120 8320
rect -120 8250 -100 8320
rect -100 8250 -80 8320
rect 10 8250 60 8320
rect 60 8250 80 8320
rect 80 8250 150 8320
rect 150 8250 170 8320
rect 170 8250 240 8320
rect 240 8250 250 8320
rect 340 8250 350 8320
rect 350 8250 420 8320
rect 420 8250 440 8320
rect 440 8250 510 8320
rect 510 8250 530 8320
rect 530 8250 580 8320
rect 670 8250 690 8320
rect 690 8250 710 8320
rect 710 8250 780 8320
rect 780 8250 800 8320
rect 800 8250 870 8320
rect 870 8250 890 8320
rect 890 8250 910 8320
rect 1000 8250 1050 8320
rect 1050 8250 1070 8320
rect 1070 8250 1140 8320
rect 1140 8250 1160 8320
rect 1160 8250 1230 8320
rect 1230 8250 1240 8320
rect 1370 8250 1380 8320
rect 1380 8250 1450 8320
rect 1450 8250 1470 8320
rect 1470 8250 1540 8320
rect 1540 8250 1560 8320
rect 1560 8250 1610 8320
rect 1700 8250 1720 8320
rect 1720 8250 1740 8320
rect 1740 8250 1810 8320
rect 1810 8250 1830 8320
rect 1830 8250 1900 8320
rect 1900 8250 1920 8320
rect 1920 8250 1940 8320
rect 2030 8250 2080 8320
rect 2080 8250 2100 8320
rect 2100 8250 2170 8320
rect 2170 8250 2190 8320
rect 2190 8250 2260 8320
rect 2260 8250 2270 8320
rect 2360 8250 2370 8320
rect 2370 8250 2440 8320
rect 2440 8250 2460 8320
rect 2460 8250 2530 8320
rect 2530 8250 2550 8320
rect 2550 8250 2600 8320
rect 2690 8250 2710 8320
rect 2710 8250 2730 8320
rect 2730 8250 2800 8320
rect 2800 8250 2820 8320
rect 2820 8250 2890 8320
rect 2890 8250 2910 8320
rect 2910 8250 2930 8320
rect 3020 8250 3070 8320
rect 3070 8250 3090 8320
rect 3090 8250 3160 8320
rect 3160 8250 3180 8320
rect 3180 8250 3250 8320
rect 3250 8250 3260 8320
rect 3350 8250 3360 8320
rect 3360 8250 3430 8320
rect 3430 8250 3450 8320
rect 3450 8250 3520 8320
rect 3520 8250 3540 8320
rect 3540 8250 3590 8320
rect 3680 8250 3700 8320
rect 3700 8250 3720 8320
rect 3720 8250 3790 8320
rect 3790 8250 3810 8320
rect 3810 8250 3880 8320
rect 3880 8250 3900 8320
rect 3900 8250 3920 8320
rect 4010 8250 4060 8320
rect 4060 8250 4080 8320
rect 4080 8250 4150 8320
rect 4150 8250 4170 8320
rect 4170 8250 4240 8320
rect 4240 8250 4250 8320
rect 4380 8250 4390 8320
rect 4390 8250 4460 8320
rect 4460 8250 4480 8320
rect 4480 8250 4550 8320
rect 4550 8250 4570 8320
rect 4570 8250 4620 8320
rect 4710 8250 4730 8320
rect 4730 8250 4750 8320
rect 4750 8250 4820 8320
rect 4820 8250 4840 8320
rect 4840 8250 4910 8320
rect 4910 8250 4930 8320
rect 4930 8250 4950 8320
rect 5040 8250 5090 8320
rect 5090 8250 5110 8320
rect 5110 8250 5180 8320
rect 5180 8250 5200 8320
rect 5200 8250 5270 8320
rect 5270 8250 5280 8320
rect 5370 8250 5380 8320
rect 5380 8250 5450 8320
rect 5450 8250 5470 8320
rect 5470 8250 5540 8320
rect 5540 8250 5560 8320
rect 5560 8250 5610 8320
rect 5700 8250 5720 8320
rect 5720 8250 5740 8320
rect 5740 8250 5810 8320
rect 5810 8250 5830 8320
rect 5830 8250 5900 8320
rect 5900 8250 5920 8320
rect 5920 8250 5940 8320
rect 6030 8250 6080 8320
rect 6080 8250 6100 8320
rect 6100 8250 6170 8320
rect 6170 8250 6190 8320
rect 6190 8250 6260 8320
rect 6260 8250 6270 8320
rect 6360 8250 6370 8320
rect 6370 8250 6440 8320
rect 6440 8250 6460 8320
rect 6460 8250 6530 8320
rect 6530 8250 6550 8320
rect 6550 8250 6600 8320
rect 6690 8250 6710 8320
rect 6710 8250 6730 8320
rect 6730 8250 6800 8320
rect 6800 8250 6820 8320
rect 6820 8250 6890 8320
rect 6890 8250 6910 8320
rect 6910 8250 6930 8320
rect 7020 8250 7070 8320
rect 7070 8250 7090 8320
rect 7090 8250 7160 8320
rect 7160 8250 7180 8320
rect 7180 8250 7250 8320
rect 7250 8250 7260 8320
rect -4650 8220 -4410 8250
rect -4320 8220 -4080 8250
rect -3990 8220 -3750 8250
rect -3660 8220 -3420 8250
rect -3330 8220 -3090 8250
rect -3000 8220 -2760 8250
rect -2670 8220 -2430 8250
rect -2340 8220 -2100 8250
rect -2010 8220 -1770 8250
rect -1640 8220 -1400 8250
rect -1310 8220 -1070 8250
rect -980 8220 -740 8250
rect -650 8220 -410 8250
rect -320 8220 -80 8250
rect 10 8220 250 8250
rect 340 8220 580 8250
rect 670 8220 910 8250
rect 1000 8220 1240 8250
rect 1370 8220 1610 8250
rect 1700 8220 1940 8250
rect 2030 8220 2270 8250
rect 2360 8220 2600 8250
rect 2690 8220 2930 8250
rect 3020 8220 3260 8250
rect 3350 8220 3590 8250
rect 3680 8220 3920 8250
rect 4010 8220 4250 8250
rect 4380 8220 4620 8250
rect 4710 8220 4950 8250
rect 5040 8220 5280 8250
rect 5370 8220 5610 8250
rect 5700 8220 5940 8250
rect 6030 8220 6270 8250
rect 6360 8220 6600 8250
rect 6690 8220 6930 8250
rect 7020 8220 7260 8250
rect 7640 8430 7650 8460
rect 7650 8430 7720 8460
rect 7720 8430 7740 8460
rect 7740 8430 7810 8460
rect 7810 8430 7830 8460
rect 7830 8430 7880 8460
rect 7970 8430 7990 8460
rect 7990 8430 8010 8460
rect 8010 8430 8080 8460
rect 8080 8430 8100 8460
rect 8100 8430 8170 8460
rect 8170 8430 8190 8460
rect 8190 8430 8210 8460
rect 8300 8430 8350 8460
rect 8350 8430 8370 8460
rect 8370 8430 8440 8460
rect 8440 8430 8460 8460
rect 8460 8430 8530 8460
rect 8530 8430 8540 8460
rect 8630 8430 8640 8460
rect 8640 8430 8710 8460
rect 8710 8430 8730 8460
rect 8730 8430 8800 8460
rect 8800 8430 8820 8460
rect 8820 8430 8870 8460
rect 8960 8430 8980 8460
rect 8980 8430 9000 8460
rect 9000 8430 9070 8460
rect 9070 8430 9090 8460
rect 9090 8430 9160 8460
rect 9160 8430 9180 8460
rect 9180 8430 9200 8460
rect 9290 8430 9340 8460
rect 9340 8430 9360 8460
rect 9360 8430 9430 8460
rect 9430 8430 9450 8460
rect 9450 8430 9520 8460
rect 9520 8430 9530 8460
rect 9620 8430 9630 8460
rect 9630 8430 9700 8460
rect 9700 8430 9720 8460
rect 9720 8430 9790 8460
rect 9790 8430 9810 8460
rect 9810 8430 9860 8460
rect 9950 8430 9970 8460
rect 9970 8430 9990 8460
rect 9990 8430 10060 8460
rect 10060 8430 10080 8460
rect 10080 8430 10150 8460
rect 10150 8430 10170 8460
rect 10170 8430 10190 8460
rect 10280 8430 10330 8460
rect 10330 8430 10350 8460
rect 10350 8430 10420 8460
rect 10420 8430 10440 8460
rect 10440 8430 10510 8460
rect 10510 8430 10520 8460
rect 10650 8430 10660 8460
rect 10660 8430 10730 8460
rect 10730 8430 10750 8460
rect 10750 8430 10820 8460
rect 10820 8430 10840 8460
rect 10840 8430 10890 8460
rect 10980 8430 11000 8460
rect 11000 8430 11020 8460
rect 11020 8430 11090 8460
rect 11090 8430 11110 8460
rect 11110 8430 11180 8460
rect 11180 8430 11200 8460
rect 11200 8430 11220 8460
rect 11310 8430 11360 8460
rect 11360 8430 11380 8460
rect 11380 8430 11450 8460
rect 11450 8430 11470 8460
rect 11470 8430 11540 8460
rect 11540 8430 11550 8460
rect 11640 8430 11650 8460
rect 11650 8430 11720 8460
rect 11720 8430 11740 8460
rect 11740 8430 11810 8460
rect 11810 8430 11830 8460
rect 11830 8430 11880 8460
rect 11970 8430 11990 8460
rect 11990 8430 12010 8460
rect 12010 8430 12080 8460
rect 12080 8430 12100 8460
rect 12100 8430 12170 8460
rect 12170 8430 12190 8460
rect 12190 8430 12210 8460
rect 12300 8430 12350 8460
rect 12350 8430 12370 8460
rect 12370 8430 12440 8460
rect 12440 8430 12460 8460
rect 12460 8430 12530 8460
rect 12530 8430 12540 8460
rect 12630 8430 12640 8460
rect 12640 8430 12710 8460
rect 12710 8430 12730 8460
rect 12730 8430 12800 8460
rect 12800 8430 12820 8460
rect 12820 8430 12870 8460
rect 12960 8430 12980 8460
rect 12980 8430 13000 8460
rect 13000 8430 13070 8460
rect 13070 8430 13090 8460
rect 13090 8430 13160 8460
rect 13160 8430 13180 8460
rect 13180 8430 13200 8460
rect 13290 8430 13340 8460
rect 13340 8430 13360 8460
rect 13360 8430 13430 8460
rect 13430 8430 13450 8460
rect 13450 8430 13520 8460
rect 13520 8430 13530 8460
rect 13660 8430 13670 8460
rect 13670 8430 13740 8460
rect 13740 8430 13760 8460
rect 13760 8430 13830 8460
rect 13830 8430 13850 8460
rect 13850 8430 13900 8460
rect 13990 8430 14010 8460
rect 14010 8430 14030 8460
rect 14030 8430 14100 8460
rect 14100 8430 14120 8460
rect 14120 8430 14190 8460
rect 14190 8430 14210 8460
rect 14210 8430 14230 8460
rect 14320 8430 14370 8460
rect 14370 8430 14390 8460
rect 14390 8430 14460 8460
rect 14460 8430 14480 8460
rect 14480 8430 14550 8460
rect 14550 8430 14560 8460
rect 14650 8430 14660 8460
rect 14660 8430 14730 8460
rect 14730 8430 14750 8460
rect 14750 8430 14820 8460
rect 14820 8430 14840 8460
rect 14840 8430 14890 8460
rect 14980 8430 15000 8460
rect 15000 8430 15020 8460
rect 15020 8430 15090 8460
rect 15090 8430 15110 8460
rect 15110 8430 15180 8460
rect 15180 8430 15200 8460
rect 15200 8430 15220 8460
rect 15310 8430 15360 8460
rect 15360 8430 15380 8460
rect 15380 8430 15450 8460
rect 15450 8430 15470 8460
rect 15470 8430 15540 8460
rect 15540 8430 15550 8460
rect 15640 8430 15650 8460
rect 15650 8430 15720 8460
rect 15720 8430 15740 8460
rect 15740 8430 15810 8460
rect 15810 8430 15830 8460
rect 15830 8430 15880 8460
rect 15970 8430 15990 8460
rect 15990 8430 16010 8460
rect 16010 8430 16080 8460
rect 16080 8430 16100 8460
rect 16100 8430 16170 8460
rect 16170 8430 16190 8460
rect 16190 8430 16210 8460
rect 16300 8430 16350 8460
rect 16350 8430 16370 8460
rect 16370 8430 16440 8460
rect 16440 8430 16460 8460
rect 16460 8430 16530 8460
rect 16530 8430 16540 8460
rect 16670 8430 16680 8460
rect 16680 8430 16750 8460
rect 16750 8430 16770 8460
rect 16770 8430 16840 8460
rect 16840 8430 16860 8460
rect 16860 8430 16910 8460
rect 17000 8430 17020 8460
rect 17020 8430 17040 8460
rect 17040 8430 17110 8460
rect 17110 8430 17130 8460
rect 17130 8430 17200 8460
rect 17200 8430 17220 8460
rect 17220 8430 17240 8460
rect 17330 8430 17380 8460
rect 17380 8430 17400 8460
rect 17400 8430 17470 8460
rect 17470 8430 17490 8460
rect 17490 8430 17560 8460
rect 17560 8430 17570 8460
rect 17660 8430 17670 8460
rect 17670 8430 17740 8460
rect 17740 8430 17760 8460
rect 17760 8430 17830 8460
rect 17830 8430 17850 8460
rect 17850 8430 17900 8460
rect 17990 8430 18010 8460
rect 18010 8430 18030 8460
rect 18030 8430 18100 8460
rect 18100 8430 18120 8460
rect 18120 8430 18190 8460
rect 18190 8430 18210 8460
rect 18210 8430 18230 8460
rect 18320 8430 18370 8460
rect 18370 8430 18390 8460
rect 18390 8430 18460 8460
rect 18460 8430 18480 8460
rect 18480 8430 18550 8460
rect 18550 8430 18560 8460
rect 18650 8430 18660 8460
rect 18660 8430 18730 8460
rect 18730 8430 18750 8460
rect 18750 8430 18820 8460
rect 18820 8430 18840 8460
rect 18840 8430 18890 8460
rect 18980 8430 19000 8460
rect 19000 8430 19020 8460
rect 19020 8430 19090 8460
rect 19090 8430 19110 8460
rect 19110 8430 19180 8460
rect 19180 8430 19200 8460
rect 19200 8430 19220 8460
rect 19310 8430 19360 8460
rect 19360 8430 19380 8460
rect 19380 8430 19450 8460
rect 19450 8430 19470 8460
rect 19470 8430 19540 8460
rect 19540 8430 19550 8460
rect 7640 8410 7880 8430
rect 7970 8410 8210 8430
rect 8300 8410 8540 8430
rect 8630 8410 8870 8430
rect 8960 8410 9200 8430
rect 9290 8410 9530 8430
rect 9620 8410 9860 8430
rect 9950 8410 10190 8430
rect 10280 8410 10520 8430
rect 10650 8410 10890 8430
rect 10980 8410 11220 8430
rect 11310 8410 11550 8430
rect 11640 8410 11880 8430
rect 11970 8410 12210 8430
rect 12300 8410 12540 8430
rect 12630 8410 12870 8430
rect 12960 8410 13200 8430
rect 13290 8410 13530 8430
rect 13660 8410 13900 8430
rect 13990 8410 14230 8430
rect 14320 8410 14560 8430
rect 14650 8410 14890 8430
rect 14980 8410 15220 8430
rect 15310 8410 15550 8430
rect 15640 8410 15880 8430
rect 15970 8410 16210 8430
rect 16300 8410 16540 8430
rect 16670 8410 16910 8430
rect 17000 8410 17240 8430
rect 17330 8410 17570 8430
rect 17660 8410 17900 8430
rect 17990 8410 18230 8430
rect 18320 8410 18560 8430
rect 18650 8410 18890 8430
rect 18980 8410 19220 8430
rect 19310 8410 19550 8430
rect 7640 8340 7650 8410
rect 7650 8340 7720 8410
rect 7720 8340 7740 8410
rect 7740 8340 7810 8410
rect 7810 8340 7830 8410
rect 7830 8340 7880 8410
rect 7970 8340 7990 8410
rect 7990 8340 8010 8410
rect 8010 8340 8080 8410
rect 8080 8340 8100 8410
rect 8100 8340 8170 8410
rect 8170 8340 8190 8410
rect 8190 8340 8210 8410
rect 8300 8340 8350 8410
rect 8350 8340 8370 8410
rect 8370 8340 8440 8410
rect 8440 8340 8460 8410
rect 8460 8340 8530 8410
rect 8530 8340 8540 8410
rect 8630 8340 8640 8410
rect 8640 8340 8710 8410
rect 8710 8340 8730 8410
rect 8730 8340 8800 8410
rect 8800 8340 8820 8410
rect 8820 8340 8870 8410
rect 8960 8340 8980 8410
rect 8980 8340 9000 8410
rect 9000 8340 9070 8410
rect 9070 8340 9090 8410
rect 9090 8340 9160 8410
rect 9160 8340 9180 8410
rect 9180 8340 9200 8410
rect 9290 8340 9340 8410
rect 9340 8340 9360 8410
rect 9360 8340 9430 8410
rect 9430 8340 9450 8410
rect 9450 8340 9520 8410
rect 9520 8340 9530 8410
rect 9620 8340 9630 8410
rect 9630 8340 9700 8410
rect 9700 8340 9720 8410
rect 9720 8340 9790 8410
rect 9790 8340 9810 8410
rect 9810 8340 9860 8410
rect 9950 8340 9970 8410
rect 9970 8340 9990 8410
rect 9990 8340 10060 8410
rect 10060 8340 10080 8410
rect 10080 8340 10150 8410
rect 10150 8340 10170 8410
rect 10170 8340 10190 8410
rect 10280 8340 10330 8410
rect 10330 8340 10350 8410
rect 10350 8340 10420 8410
rect 10420 8340 10440 8410
rect 10440 8340 10510 8410
rect 10510 8340 10520 8410
rect 10650 8340 10660 8410
rect 10660 8340 10730 8410
rect 10730 8340 10750 8410
rect 10750 8340 10820 8410
rect 10820 8340 10840 8410
rect 10840 8340 10890 8410
rect 10980 8340 11000 8410
rect 11000 8340 11020 8410
rect 11020 8340 11090 8410
rect 11090 8340 11110 8410
rect 11110 8340 11180 8410
rect 11180 8340 11200 8410
rect 11200 8340 11220 8410
rect 11310 8340 11360 8410
rect 11360 8340 11380 8410
rect 11380 8340 11450 8410
rect 11450 8340 11470 8410
rect 11470 8340 11540 8410
rect 11540 8340 11550 8410
rect 11640 8340 11650 8410
rect 11650 8340 11720 8410
rect 11720 8340 11740 8410
rect 11740 8340 11810 8410
rect 11810 8340 11830 8410
rect 11830 8340 11880 8410
rect 11970 8340 11990 8410
rect 11990 8340 12010 8410
rect 12010 8340 12080 8410
rect 12080 8340 12100 8410
rect 12100 8340 12170 8410
rect 12170 8340 12190 8410
rect 12190 8340 12210 8410
rect 12300 8340 12350 8410
rect 12350 8340 12370 8410
rect 12370 8340 12440 8410
rect 12440 8340 12460 8410
rect 12460 8340 12530 8410
rect 12530 8340 12540 8410
rect 12630 8340 12640 8410
rect 12640 8340 12710 8410
rect 12710 8340 12730 8410
rect 12730 8340 12800 8410
rect 12800 8340 12820 8410
rect 12820 8340 12870 8410
rect 12960 8340 12980 8410
rect 12980 8340 13000 8410
rect 13000 8340 13070 8410
rect 13070 8340 13090 8410
rect 13090 8340 13160 8410
rect 13160 8340 13180 8410
rect 13180 8340 13200 8410
rect 13290 8340 13340 8410
rect 13340 8340 13360 8410
rect 13360 8340 13430 8410
rect 13430 8340 13450 8410
rect 13450 8340 13520 8410
rect 13520 8340 13530 8410
rect 13660 8340 13670 8410
rect 13670 8340 13740 8410
rect 13740 8340 13760 8410
rect 13760 8340 13830 8410
rect 13830 8340 13850 8410
rect 13850 8340 13900 8410
rect 13990 8340 14010 8410
rect 14010 8340 14030 8410
rect 14030 8340 14100 8410
rect 14100 8340 14120 8410
rect 14120 8340 14190 8410
rect 14190 8340 14210 8410
rect 14210 8340 14230 8410
rect 14320 8340 14370 8410
rect 14370 8340 14390 8410
rect 14390 8340 14460 8410
rect 14460 8340 14480 8410
rect 14480 8340 14550 8410
rect 14550 8340 14560 8410
rect 14650 8340 14660 8410
rect 14660 8340 14730 8410
rect 14730 8340 14750 8410
rect 14750 8340 14820 8410
rect 14820 8340 14840 8410
rect 14840 8340 14890 8410
rect 14980 8340 15000 8410
rect 15000 8340 15020 8410
rect 15020 8340 15090 8410
rect 15090 8340 15110 8410
rect 15110 8340 15180 8410
rect 15180 8340 15200 8410
rect 15200 8340 15220 8410
rect 15310 8340 15360 8410
rect 15360 8340 15380 8410
rect 15380 8340 15450 8410
rect 15450 8340 15470 8410
rect 15470 8340 15540 8410
rect 15540 8340 15550 8410
rect 15640 8340 15650 8410
rect 15650 8340 15720 8410
rect 15720 8340 15740 8410
rect 15740 8340 15810 8410
rect 15810 8340 15830 8410
rect 15830 8340 15880 8410
rect 15970 8340 15990 8410
rect 15990 8340 16010 8410
rect 16010 8340 16080 8410
rect 16080 8340 16100 8410
rect 16100 8340 16170 8410
rect 16170 8340 16190 8410
rect 16190 8340 16210 8410
rect 16300 8340 16350 8410
rect 16350 8340 16370 8410
rect 16370 8340 16440 8410
rect 16440 8340 16460 8410
rect 16460 8340 16530 8410
rect 16530 8340 16540 8410
rect 16670 8340 16680 8410
rect 16680 8340 16750 8410
rect 16750 8340 16770 8410
rect 16770 8340 16840 8410
rect 16840 8340 16860 8410
rect 16860 8340 16910 8410
rect 17000 8340 17020 8410
rect 17020 8340 17040 8410
rect 17040 8340 17110 8410
rect 17110 8340 17130 8410
rect 17130 8340 17200 8410
rect 17200 8340 17220 8410
rect 17220 8340 17240 8410
rect 17330 8340 17380 8410
rect 17380 8340 17400 8410
rect 17400 8340 17470 8410
rect 17470 8340 17490 8410
rect 17490 8340 17560 8410
rect 17560 8340 17570 8410
rect 17660 8340 17670 8410
rect 17670 8340 17740 8410
rect 17740 8340 17760 8410
rect 17760 8340 17830 8410
rect 17830 8340 17850 8410
rect 17850 8340 17900 8410
rect 17990 8340 18010 8410
rect 18010 8340 18030 8410
rect 18030 8340 18100 8410
rect 18100 8340 18120 8410
rect 18120 8340 18190 8410
rect 18190 8340 18210 8410
rect 18210 8340 18230 8410
rect 18320 8340 18370 8410
rect 18370 8340 18390 8410
rect 18390 8340 18460 8410
rect 18460 8340 18480 8410
rect 18480 8340 18550 8410
rect 18550 8340 18560 8410
rect 18650 8340 18660 8410
rect 18660 8340 18730 8410
rect 18730 8340 18750 8410
rect 18750 8340 18820 8410
rect 18820 8340 18840 8410
rect 18840 8340 18890 8410
rect 18980 8340 19000 8410
rect 19000 8340 19020 8410
rect 19020 8340 19090 8410
rect 19090 8340 19110 8410
rect 19110 8340 19180 8410
rect 19180 8340 19200 8410
rect 19200 8340 19220 8410
rect 19310 8340 19360 8410
rect 19360 8340 19380 8410
rect 19380 8340 19450 8410
rect 19450 8340 19470 8410
rect 19470 8340 19540 8410
rect 19540 8340 19550 8410
rect 7640 8320 7880 8340
rect 7970 8320 8210 8340
rect 8300 8320 8540 8340
rect 8630 8320 8870 8340
rect 8960 8320 9200 8340
rect 9290 8320 9530 8340
rect 9620 8320 9860 8340
rect 9950 8320 10190 8340
rect 10280 8320 10520 8340
rect 10650 8320 10890 8340
rect 10980 8320 11220 8340
rect 11310 8320 11550 8340
rect 11640 8320 11880 8340
rect 11970 8320 12210 8340
rect 12300 8320 12540 8340
rect 12630 8320 12870 8340
rect 12960 8320 13200 8340
rect 13290 8320 13530 8340
rect 13660 8320 13900 8340
rect 13990 8320 14230 8340
rect 14320 8320 14560 8340
rect 14650 8320 14890 8340
rect 14980 8320 15220 8340
rect 15310 8320 15550 8340
rect 15640 8320 15880 8340
rect 15970 8320 16210 8340
rect 16300 8320 16540 8340
rect 16670 8320 16910 8340
rect 17000 8320 17240 8340
rect 17330 8320 17570 8340
rect 17660 8320 17900 8340
rect 17990 8320 18230 8340
rect 18320 8320 18560 8340
rect 18650 8320 18890 8340
rect 18980 8320 19220 8340
rect 19310 8320 19550 8340
rect 7640 8250 7650 8320
rect 7650 8250 7720 8320
rect 7720 8250 7740 8320
rect 7740 8250 7810 8320
rect 7810 8250 7830 8320
rect 7830 8250 7880 8320
rect 7970 8250 7990 8320
rect 7990 8250 8010 8320
rect 8010 8250 8080 8320
rect 8080 8250 8100 8320
rect 8100 8250 8170 8320
rect 8170 8250 8190 8320
rect 8190 8250 8210 8320
rect 8300 8250 8350 8320
rect 8350 8250 8370 8320
rect 8370 8250 8440 8320
rect 8440 8250 8460 8320
rect 8460 8250 8530 8320
rect 8530 8250 8540 8320
rect 8630 8250 8640 8320
rect 8640 8250 8710 8320
rect 8710 8250 8730 8320
rect 8730 8250 8800 8320
rect 8800 8250 8820 8320
rect 8820 8250 8870 8320
rect 8960 8250 8980 8320
rect 8980 8250 9000 8320
rect 9000 8250 9070 8320
rect 9070 8250 9090 8320
rect 9090 8250 9160 8320
rect 9160 8250 9180 8320
rect 9180 8250 9200 8320
rect 9290 8250 9340 8320
rect 9340 8250 9360 8320
rect 9360 8250 9430 8320
rect 9430 8250 9450 8320
rect 9450 8250 9520 8320
rect 9520 8250 9530 8320
rect 9620 8250 9630 8320
rect 9630 8250 9700 8320
rect 9700 8250 9720 8320
rect 9720 8250 9790 8320
rect 9790 8250 9810 8320
rect 9810 8250 9860 8320
rect 9950 8250 9970 8320
rect 9970 8250 9990 8320
rect 9990 8250 10060 8320
rect 10060 8250 10080 8320
rect 10080 8250 10150 8320
rect 10150 8250 10170 8320
rect 10170 8250 10190 8320
rect 10280 8250 10330 8320
rect 10330 8250 10350 8320
rect 10350 8250 10420 8320
rect 10420 8250 10440 8320
rect 10440 8250 10510 8320
rect 10510 8250 10520 8320
rect 10650 8250 10660 8320
rect 10660 8250 10730 8320
rect 10730 8250 10750 8320
rect 10750 8250 10820 8320
rect 10820 8250 10840 8320
rect 10840 8250 10890 8320
rect 10980 8250 11000 8320
rect 11000 8250 11020 8320
rect 11020 8250 11090 8320
rect 11090 8250 11110 8320
rect 11110 8250 11180 8320
rect 11180 8250 11200 8320
rect 11200 8250 11220 8320
rect 11310 8250 11360 8320
rect 11360 8250 11380 8320
rect 11380 8250 11450 8320
rect 11450 8250 11470 8320
rect 11470 8250 11540 8320
rect 11540 8250 11550 8320
rect 11640 8250 11650 8320
rect 11650 8250 11720 8320
rect 11720 8250 11740 8320
rect 11740 8250 11810 8320
rect 11810 8250 11830 8320
rect 11830 8250 11880 8320
rect 11970 8250 11990 8320
rect 11990 8250 12010 8320
rect 12010 8250 12080 8320
rect 12080 8250 12100 8320
rect 12100 8250 12170 8320
rect 12170 8250 12190 8320
rect 12190 8250 12210 8320
rect 12300 8250 12350 8320
rect 12350 8250 12370 8320
rect 12370 8250 12440 8320
rect 12440 8250 12460 8320
rect 12460 8250 12530 8320
rect 12530 8250 12540 8320
rect 12630 8250 12640 8320
rect 12640 8250 12710 8320
rect 12710 8250 12730 8320
rect 12730 8250 12800 8320
rect 12800 8250 12820 8320
rect 12820 8250 12870 8320
rect 12960 8250 12980 8320
rect 12980 8250 13000 8320
rect 13000 8250 13070 8320
rect 13070 8250 13090 8320
rect 13090 8250 13160 8320
rect 13160 8250 13180 8320
rect 13180 8250 13200 8320
rect 13290 8250 13340 8320
rect 13340 8250 13360 8320
rect 13360 8250 13430 8320
rect 13430 8250 13450 8320
rect 13450 8250 13520 8320
rect 13520 8250 13530 8320
rect 13660 8250 13670 8320
rect 13670 8250 13740 8320
rect 13740 8250 13760 8320
rect 13760 8250 13830 8320
rect 13830 8250 13850 8320
rect 13850 8250 13900 8320
rect 13990 8250 14010 8320
rect 14010 8250 14030 8320
rect 14030 8250 14100 8320
rect 14100 8250 14120 8320
rect 14120 8250 14190 8320
rect 14190 8250 14210 8320
rect 14210 8250 14230 8320
rect 14320 8250 14370 8320
rect 14370 8250 14390 8320
rect 14390 8250 14460 8320
rect 14460 8250 14480 8320
rect 14480 8250 14550 8320
rect 14550 8250 14560 8320
rect 14650 8250 14660 8320
rect 14660 8250 14730 8320
rect 14730 8250 14750 8320
rect 14750 8250 14820 8320
rect 14820 8250 14840 8320
rect 14840 8250 14890 8320
rect 14980 8250 15000 8320
rect 15000 8250 15020 8320
rect 15020 8250 15090 8320
rect 15090 8250 15110 8320
rect 15110 8250 15180 8320
rect 15180 8250 15200 8320
rect 15200 8250 15220 8320
rect 15310 8250 15360 8320
rect 15360 8250 15380 8320
rect 15380 8250 15450 8320
rect 15450 8250 15470 8320
rect 15470 8250 15540 8320
rect 15540 8250 15550 8320
rect 15640 8250 15650 8320
rect 15650 8250 15720 8320
rect 15720 8250 15740 8320
rect 15740 8250 15810 8320
rect 15810 8250 15830 8320
rect 15830 8250 15880 8320
rect 15970 8250 15990 8320
rect 15990 8250 16010 8320
rect 16010 8250 16080 8320
rect 16080 8250 16100 8320
rect 16100 8250 16170 8320
rect 16170 8250 16190 8320
rect 16190 8250 16210 8320
rect 16300 8250 16350 8320
rect 16350 8250 16370 8320
rect 16370 8250 16440 8320
rect 16440 8250 16460 8320
rect 16460 8250 16530 8320
rect 16530 8250 16540 8320
rect 16670 8250 16680 8320
rect 16680 8250 16750 8320
rect 16750 8250 16770 8320
rect 16770 8250 16840 8320
rect 16840 8250 16860 8320
rect 16860 8250 16910 8320
rect 17000 8250 17020 8320
rect 17020 8250 17040 8320
rect 17040 8250 17110 8320
rect 17110 8250 17130 8320
rect 17130 8250 17200 8320
rect 17200 8250 17220 8320
rect 17220 8250 17240 8320
rect 17330 8250 17380 8320
rect 17380 8250 17400 8320
rect 17400 8250 17470 8320
rect 17470 8250 17490 8320
rect 17490 8250 17560 8320
rect 17560 8250 17570 8320
rect 17660 8250 17670 8320
rect 17670 8250 17740 8320
rect 17740 8250 17760 8320
rect 17760 8250 17830 8320
rect 17830 8250 17850 8320
rect 17850 8250 17900 8320
rect 17990 8250 18010 8320
rect 18010 8250 18030 8320
rect 18030 8250 18100 8320
rect 18100 8250 18120 8320
rect 18120 8250 18190 8320
rect 18190 8250 18210 8320
rect 18210 8250 18230 8320
rect 18320 8250 18370 8320
rect 18370 8250 18390 8320
rect 18390 8250 18460 8320
rect 18460 8250 18480 8320
rect 18480 8250 18550 8320
rect 18550 8250 18560 8320
rect 18650 8250 18660 8320
rect 18660 8250 18730 8320
rect 18730 8250 18750 8320
rect 18750 8250 18820 8320
rect 18820 8250 18840 8320
rect 18840 8250 18890 8320
rect 18980 8250 19000 8320
rect 19000 8250 19020 8320
rect 19020 8250 19090 8320
rect 19090 8250 19110 8320
rect 19110 8250 19180 8320
rect 19180 8250 19200 8320
rect 19200 8250 19220 8320
rect 19310 8250 19360 8320
rect 19360 8250 19380 8320
rect 19380 8250 19450 8320
rect 19450 8250 19470 8320
rect 19470 8250 19540 8320
rect 19540 8250 19550 8320
rect 7640 8220 7880 8250
rect 7970 8220 8210 8250
rect 8300 8220 8540 8250
rect 8630 8220 8870 8250
rect 8960 8220 9200 8250
rect 9290 8220 9530 8250
rect 9620 8220 9860 8250
rect 9950 8220 10190 8250
rect 10280 8220 10520 8250
rect 10650 8220 10890 8250
rect 10980 8220 11220 8250
rect 11310 8220 11550 8250
rect 11640 8220 11880 8250
rect 11970 8220 12210 8250
rect 12300 8220 12540 8250
rect 12630 8220 12870 8250
rect 12960 8220 13200 8250
rect 13290 8220 13530 8250
rect 13660 8220 13900 8250
rect 13990 8220 14230 8250
rect 14320 8220 14560 8250
rect 14650 8220 14890 8250
rect 14980 8220 15220 8250
rect 15310 8220 15550 8250
rect 15640 8220 15880 8250
rect 15970 8220 16210 8250
rect 16300 8220 16540 8250
rect 16670 8220 16910 8250
rect 17000 8220 17240 8250
rect 17330 8220 17570 8250
rect 17660 8220 17900 8250
rect 17990 8220 18230 8250
rect 18320 8220 18560 8250
rect 18650 8220 18890 8250
rect 18980 8220 19220 8250
rect 19310 8220 19550 8250
rect 21110 7210 21480 7270
rect 21110 7140 21160 7210
rect 21160 7140 21200 7210
rect 21200 7140 21270 7210
rect 21270 7140 21310 7210
rect 21310 7140 21380 7210
rect 21380 7140 21420 7210
rect 21420 7140 21480 7210
rect 21110 7100 21480 7140
rect 21110 7030 21160 7100
rect 21160 7030 21200 7100
rect 21200 7030 21270 7100
rect 21270 7030 21310 7100
rect 21310 7030 21380 7100
rect 21380 7030 21420 7100
rect 21420 7030 21480 7100
rect 23510 7210 23880 7270
rect 23510 7140 23560 7210
rect 23560 7140 23600 7210
rect 23600 7140 23670 7210
rect 23670 7140 23710 7210
rect 23710 7140 23780 7210
rect 23780 7140 23820 7210
rect 23820 7140 23880 7210
rect 23510 7100 23880 7140
rect 23510 7030 23560 7100
rect 23560 7030 23600 7100
rect 23600 7030 23670 7100
rect 23670 7030 23710 7100
rect 23710 7030 23780 7100
rect 23780 7030 23820 7100
rect 23820 7030 23880 7100
rect 1720 6850 1960 6910
rect 2050 6850 2290 6910
rect 2390 6850 2630 6910
rect 2720 6850 2960 6910
rect 1720 6780 1750 6850
rect 1750 6780 1790 6850
rect 1790 6780 1860 6850
rect 1860 6780 1900 6850
rect 1900 6780 1960 6850
rect 2050 6780 2080 6850
rect 2080 6780 2120 6850
rect 2120 6780 2190 6850
rect 2190 6780 2230 6850
rect 2230 6780 2290 6850
rect 2390 6780 2410 6850
rect 2410 6780 2450 6850
rect 2450 6780 2520 6850
rect 2520 6780 2560 6850
rect 2560 6780 2630 6850
rect 2720 6780 2740 6850
rect 2740 6780 2780 6850
rect 2780 6780 2850 6850
rect 2850 6780 2890 6850
rect 2890 6780 2960 6850
rect 1720 6740 1960 6780
rect 2050 6740 2290 6780
rect 2390 6740 2630 6780
rect 2720 6740 2960 6780
rect 1720 6670 1750 6740
rect 1750 6670 1790 6740
rect 1790 6670 1860 6740
rect 1860 6670 1900 6740
rect 1900 6670 1960 6740
rect 2050 6670 2080 6740
rect 2080 6670 2120 6740
rect 2120 6670 2190 6740
rect 2190 6670 2230 6740
rect 2230 6670 2290 6740
rect 2390 6670 2410 6740
rect 2410 6670 2450 6740
rect 2450 6670 2520 6740
rect 2520 6670 2560 6740
rect 2560 6670 2630 6740
rect 2720 6670 2740 6740
rect 2740 6670 2780 6740
rect 2780 6670 2850 6740
rect 2850 6670 2890 6740
rect 2890 6670 2960 6740
rect 11940 6880 12180 6940
rect 12270 6880 12510 6940
rect 12610 6880 12850 6940
rect 12940 6880 13180 6940
rect 11940 6810 11970 6880
rect 11970 6810 12010 6880
rect 12010 6810 12080 6880
rect 12080 6810 12120 6880
rect 12120 6810 12180 6880
rect 12270 6810 12300 6880
rect 12300 6810 12340 6880
rect 12340 6810 12410 6880
rect 12410 6810 12450 6880
rect 12450 6810 12510 6880
rect 12610 6810 12630 6880
rect 12630 6810 12670 6880
rect 12670 6810 12740 6880
rect 12740 6810 12780 6880
rect 12780 6810 12850 6880
rect 12940 6810 12960 6880
rect 12960 6810 13000 6880
rect 13000 6810 13070 6880
rect 13070 6810 13110 6880
rect 13110 6810 13180 6880
rect 11940 6770 12180 6810
rect 12270 6770 12510 6810
rect 12610 6770 12850 6810
rect 12940 6770 13180 6810
rect 11940 6700 11970 6770
rect 11970 6700 12010 6770
rect 12010 6700 12080 6770
rect 12080 6700 12120 6770
rect 12120 6700 12180 6770
rect 12270 6700 12300 6770
rect 12300 6700 12340 6770
rect 12340 6700 12410 6770
rect 12410 6700 12450 6770
rect 12450 6700 12510 6770
rect 12610 6700 12630 6770
rect 12630 6700 12670 6770
rect 12670 6700 12740 6770
rect 12740 6700 12780 6770
rect 12780 6700 12850 6770
rect 12940 6700 12960 6770
rect 12960 6700 13000 6770
rect 13000 6700 13070 6770
rect 13070 6700 13110 6770
rect 13110 6700 13180 6770
rect 20080 2530 20140 2600
rect 20140 2530 20180 2600
rect 20180 2530 20250 2600
rect 20250 2530 20290 2600
rect 20290 2530 20360 2600
rect 20360 2530 20400 2600
rect 20400 2530 20450 2600
rect 20080 2490 20450 2530
rect 20080 2420 20140 2490
rect 20140 2420 20180 2490
rect 20180 2420 20250 2490
rect 20250 2420 20290 2490
rect 20290 2420 20360 2490
rect 20360 2420 20400 2490
rect 20400 2420 20450 2490
rect 20080 2360 20450 2420
rect 24560 2530 24620 2600
rect 24620 2530 24660 2600
rect 24660 2530 24730 2600
rect 24730 2530 24770 2600
rect 24770 2530 24840 2600
rect 24840 2530 24880 2600
rect 24880 2530 24930 2600
rect 24560 2490 24930 2530
rect 24560 2420 24620 2490
rect 24620 2420 24660 2490
rect 24660 2420 24730 2490
rect 24730 2420 24770 2490
rect 24770 2420 24840 2490
rect 24840 2420 24880 2490
rect 24880 2420 24930 2490
rect 24560 2360 24930 2420
rect 1260 -860 1330 -790
rect 1330 -860 1370 -790
rect 1370 -860 1440 -790
rect 1440 -860 1480 -790
rect 1480 -860 1500 -790
rect 1590 -860 1660 -790
rect 1660 -860 1700 -790
rect 1700 -860 1770 -790
rect 1770 -860 1810 -790
rect 1810 -860 1830 -790
rect 1930 -860 1990 -790
rect 1990 -860 2030 -790
rect 2030 -860 2100 -790
rect 2100 -860 2140 -790
rect 2140 -860 2170 -790
rect 2260 -860 2320 -790
rect 2320 -860 2360 -790
rect 2360 -860 2430 -790
rect 2430 -860 2470 -790
rect 2470 -860 2500 -790
rect 1260 -900 1500 -860
rect 1590 -900 1830 -860
rect 1930 -900 2170 -860
rect 2260 -900 2500 -860
rect 1260 -970 1330 -900
rect 1330 -970 1370 -900
rect 1370 -970 1440 -900
rect 1440 -970 1480 -900
rect 1480 -970 1500 -900
rect 1590 -970 1660 -900
rect 1660 -970 1700 -900
rect 1700 -970 1770 -900
rect 1770 -970 1810 -900
rect 1810 -970 1830 -900
rect 1930 -970 1990 -900
rect 1990 -970 2030 -900
rect 2030 -970 2100 -900
rect 2100 -970 2140 -900
rect 2140 -970 2170 -900
rect 2260 -970 2320 -900
rect 2320 -970 2360 -900
rect 2360 -970 2430 -900
rect 2430 -970 2470 -900
rect 2470 -970 2500 -900
rect 1260 -1030 1500 -970
rect 1590 -1030 1830 -970
rect 1930 -1030 2170 -970
rect 2260 -1030 2500 -970
rect 12400 -860 12430 -790
rect 12430 -860 12470 -790
rect 12470 -860 12540 -790
rect 12540 -860 12580 -790
rect 12580 -860 12640 -790
rect 12730 -860 12760 -790
rect 12760 -860 12800 -790
rect 12800 -860 12870 -790
rect 12870 -860 12910 -790
rect 12910 -860 12970 -790
rect 13070 -860 13090 -790
rect 13090 -860 13130 -790
rect 13130 -860 13200 -790
rect 13200 -860 13240 -790
rect 13240 -860 13310 -790
rect 13400 -860 13420 -790
rect 13420 -860 13460 -790
rect 13460 -860 13530 -790
rect 13530 -860 13570 -790
rect 13570 -860 13640 -790
rect 12400 -900 12640 -860
rect 12730 -900 12970 -860
rect 13070 -900 13310 -860
rect 13400 -900 13640 -860
rect 12400 -970 12430 -900
rect 12430 -970 12470 -900
rect 12470 -970 12540 -900
rect 12540 -970 12580 -900
rect 12580 -970 12640 -900
rect 12730 -970 12760 -900
rect 12760 -970 12800 -900
rect 12800 -970 12870 -900
rect 12870 -970 12910 -900
rect 12910 -970 12970 -900
rect 13070 -970 13090 -900
rect 13090 -970 13130 -900
rect 13130 -970 13200 -900
rect 13200 -970 13240 -900
rect 13240 -970 13310 -900
rect 13400 -970 13420 -900
rect 13420 -970 13460 -900
rect 13460 -970 13530 -900
rect 13530 -970 13570 -900
rect 13570 -970 13640 -900
rect 12400 -1030 12640 -970
rect 12730 -1030 12970 -970
rect 13070 -1030 13310 -970
rect 13400 -1030 13640 -970
rect 1720 -2780 1960 -2720
rect 2050 -2780 2290 -2720
rect 2390 -2780 2630 -2720
rect 2720 -2780 2960 -2720
rect 1720 -2850 1750 -2780
rect 1750 -2850 1790 -2780
rect 1790 -2850 1860 -2780
rect 1860 -2850 1900 -2780
rect 1900 -2850 1960 -2780
rect 2050 -2850 2080 -2780
rect 2080 -2850 2120 -2780
rect 2120 -2850 2190 -2780
rect 2190 -2850 2230 -2780
rect 2230 -2850 2290 -2780
rect 2390 -2850 2410 -2780
rect 2410 -2850 2450 -2780
rect 2450 -2850 2520 -2780
rect 2520 -2850 2560 -2780
rect 2560 -2850 2630 -2780
rect 2720 -2850 2740 -2780
rect 2740 -2850 2780 -2780
rect 2780 -2850 2850 -2780
rect 2850 -2850 2890 -2780
rect 2890 -2850 2960 -2780
rect 1720 -2890 1960 -2850
rect 2050 -2890 2290 -2850
rect 2390 -2890 2630 -2850
rect 2720 -2890 2960 -2850
rect 1720 -2960 1750 -2890
rect 1750 -2960 1790 -2890
rect 1790 -2960 1860 -2890
rect 1860 -2960 1900 -2890
rect 1900 -2960 1960 -2890
rect 2050 -2960 2080 -2890
rect 2080 -2960 2120 -2890
rect 2120 -2960 2190 -2890
rect 2190 -2960 2230 -2890
rect 2230 -2960 2290 -2890
rect 2390 -2960 2410 -2890
rect 2410 -2960 2450 -2890
rect 2450 -2960 2520 -2890
rect 2520 -2960 2560 -2890
rect 2560 -2960 2630 -2890
rect 2720 -2960 2740 -2890
rect 2740 -2960 2780 -2890
rect 2780 -2960 2850 -2890
rect 2850 -2960 2890 -2890
rect 2890 -2960 2960 -2890
rect 11940 -2780 12180 -2720
rect 12270 -2780 12510 -2720
rect 12610 -2780 12850 -2720
rect 12940 -2780 13180 -2720
rect 11940 -2850 11970 -2780
rect 11970 -2850 12010 -2780
rect 12010 -2850 12080 -2780
rect 12080 -2850 12120 -2780
rect 12120 -2850 12180 -2780
rect 12270 -2850 12300 -2780
rect 12300 -2850 12340 -2780
rect 12340 -2850 12410 -2780
rect 12410 -2850 12450 -2780
rect 12450 -2850 12510 -2780
rect 12610 -2850 12630 -2780
rect 12630 -2850 12670 -2780
rect 12670 -2850 12740 -2780
rect 12740 -2850 12780 -2780
rect 12780 -2850 12850 -2780
rect 12940 -2850 12960 -2780
rect 12960 -2850 13000 -2780
rect 13000 -2850 13070 -2780
rect 13070 -2850 13110 -2780
rect 13110 -2850 13180 -2780
rect 11940 -2890 12180 -2850
rect 12270 -2890 12510 -2850
rect 12610 -2890 12850 -2850
rect 12940 -2890 13180 -2850
rect 11940 -2960 11970 -2890
rect 11970 -2960 12010 -2890
rect 12010 -2960 12080 -2890
rect 12080 -2960 12120 -2890
rect 12120 -2960 12180 -2890
rect 12270 -2960 12300 -2890
rect 12300 -2960 12340 -2890
rect 12340 -2960 12410 -2890
rect 12410 -2960 12450 -2890
rect 12450 -2960 12510 -2890
rect 12610 -2960 12630 -2890
rect 12630 -2960 12670 -2890
rect 12670 -2960 12740 -2890
rect 12740 -2960 12780 -2890
rect 12780 -2960 12850 -2890
rect 12940 -2960 12960 -2890
rect 12960 -2960 13000 -2890
rect 13000 -2960 13070 -2890
rect 13070 -2960 13110 -2890
rect 13110 -2960 13180 -2890
rect -120 -4300 -90 -4250
rect -90 -4300 -70 -4250
rect -70 -4300 0 -4250
rect 0 -4300 20 -4250
rect 20 -4300 90 -4250
rect 90 -4300 120 -4250
rect -120 -4320 120 -4300
rect -120 -4390 -90 -4320
rect -90 -4390 -70 -4320
rect -70 -4390 0 -4320
rect 0 -4390 20 -4320
rect 20 -4390 90 -4320
rect 90 -4390 120 -4320
rect -120 -4410 120 -4390
rect -120 -4480 -90 -4410
rect -90 -4480 -70 -4410
rect -70 -4480 0 -4410
rect 0 -4480 20 -4410
rect 20 -4480 90 -4410
rect 90 -4480 120 -4410
rect -120 -4490 120 -4480
rect -120 -4590 120 -4580
rect -120 -4660 -90 -4590
rect -90 -4660 -70 -4590
rect -70 -4660 0 -4590
rect 0 -4660 20 -4590
rect 20 -4660 90 -4590
rect 90 -4660 120 -4590
rect -120 -4680 120 -4660
rect -120 -4750 -90 -4680
rect -90 -4750 -70 -4680
rect -70 -4750 0 -4680
rect 0 -4750 20 -4680
rect 20 -4750 90 -4680
rect 90 -4750 120 -4680
rect -120 -4770 120 -4750
rect -120 -4820 -90 -4770
rect -90 -4820 -70 -4770
rect -70 -4820 0 -4770
rect 0 -4820 20 -4770
rect 20 -4820 90 -4770
rect 90 -4820 120 -4770
rect -120 -4930 -90 -4910
rect -90 -4930 -70 -4910
rect -70 -4930 0 -4910
rect 0 -4930 20 -4910
rect 20 -4930 90 -4910
rect 90 -4930 120 -4910
rect -120 -4950 120 -4930
rect -120 -5020 -90 -4950
rect -90 -5020 -70 -4950
rect -70 -5020 0 -4950
rect 0 -5020 20 -4950
rect 20 -5020 90 -4950
rect 90 -5020 120 -4950
rect -120 -5040 120 -5020
rect -120 -5110 -90 -5040
rect -90 -5110 -70 -5040
rect -70 -5110 0 -5040
rect 0 -5110 20 -5040
rect 20 -5110 90 -5040
rect 90 -5110 120 -5040
rect -120 -5130 120 -5110
rect -120 -5150 -90 -5130
rect -90 -5150 -70 -5130
rect -70 -5150 0 -5130
rect 0 -5150 20 -5130
rect 20 -5150 90 -5130
rect 90 -5150 120 -5130
rect -120 -5290 -90 -5240
rect -90 -5290 -70 -5240
rect -70 -5290 0 -5240
rect 0 -5290 20 -5240
rect 20 -5290 90 -5240
rect 90 -5290 120 -5240
rect -120 -5310 120 -5290
rect -120 -5380 -90 -5310
rect -90 -5380 -70 -5310
rect -70 -5380 0 -5310
rect 0 -5380 20 -5310
rect 20 -5380 90 -5310
rect 90 -5380 120 -5310
rect -120 -5400 120 -5380
rect -120 -5470 -90 -5400
rect -90 -5470 -70 -5400
rect -70 -5470 0 -5400
rect 0 -5470 20 -5400
rect 20 -5470 90 -5400
rect 90 -5470 120 -5400
rect -120 -5480 120 -5470
rect 21110 920 21480 980
rect 21110 850 21160 920
rect 21160 850 21200 920
rect 21200 850 21270 920
rect 21270 850 21310 920
rect 21310 850 21380 920
rect 21380 850 21420 920
rect 21420 850 21480 920
rect 21110 810 21480 850
rect 21110 740 21160 810
rect 21160 740 21200 810
rect 21200 740 21270 810
rect 21270 740 21310 810
rect 21310 740 21380 810
rect 21380 740 21420 810
rect 21420 740 21480 810
rect 23510 920 23880 980
rect 23510 850 23560 920
rect 23560 850 23600 920
rect 23600 850 23670 920
rect 23670 850 23710 920
rect 23710 850 23780 920
rect 23780 850 23820 920
rect 23820 850 23880 920
rect 23510 810 23880 850
rect 23510 740 23560 810
rect 23560 740 23600 810
rect 23600 740 23670 810
rect 23670 740 23710 810
rect 23710 740 23780 810
rect 23780 740 23820 810
rect 23820 740 23880 810
rect 35830 7750 35860 7770
rect 35860 7750 35880 7770
rect 35880 7750 35950 7770
rect 35950 7750 35970 7770
rect 35970 7750 36040 7770
rect 36040 7750 36070 7770
rect 35830 7730 36070 7750
rect 35830 7660 35860 7730
rect 35860 7660 35880 7730
rect 35880 7660 35950 7730
rect 35950 7660 35970 7730
rect 35970 7660 36040 7730
rect 36040 7660 36070 7730
rect 35830 7640 36070 7660
rect 35830 7570 35860 7640
rect 35860 7570 35880 7640
rect 35880 7570 35950 7640
rect 35950 7570 35970 7640
rect 35970 7570 36040 7640
rect 36040 7570 36070 7640
rect 35830 7550 36070 7570
rect 35830 7530 35860 7550
rect 35860 7530 35880 7550
rect 35880 7530 35950 7550
rect 35950 7530 35970 7550
rect 35970 7530 36040 7550
rect 36040 7530 36070 7550
rect 35830 7390 35860 7440
rect 35860 7390 35880 7440
rect 35880 7390 35950 7440
rect 35950 7390 35970 7440
rect 35970 7390 36040 7440
rect 36040 7390 36070 7440
rect 35830 7370 36070 7390
rect 35830 7300 35860 7370
rect 35860 7300 35880 7370
rect 35880 7300 35950 7370
rect 35950 7300 35970 7370
rect 35970 7300 36040 7370
rect 36040 7300 36070 7370
rect 35830 7280 36070 7300
rect 35830 7210 35860 7280
rect 35860 7210 35880 7280
rect 35880 7210 35950 7280
rect 35950 7210 35970 7280
rect 35970 7210 36040 7280
rect 36040 7210 36070 7280
rect 35830 7200 36070 7210
rect 35830 7060 36070 7070
rect 35830 6990 35860 7060
rect 35860 6990 35880 7060
rect 35880 6990 35950 7060
rect 35950 6990 35970 7060
rect 35970 6990 36040 7060
rect 36040 6990 36070 7060
rect 35830 6970 36070 6990
rect 35830 6900 35860 6970
rect 35860 6900 35880 6970
rect 35880 6900 35950 6970
rect 35950 6900 35970 6970
rect 35970 6900 36040 6970
rect 36040 6900 36070 6970
rect 35830 6880 36070 6900
rect 35830 6830 35860 6880
rect 35860 6830 35880 6880
rect 35880 6830 35950 6880
rect 35950 6830 35970 6880
rect 35970 6830 36040 6880
rect 36040 6830 36070 6880
rect 35830 6720 35860 6740
rect 35860 6720 35880 6740
rect 35880 6720 35950 6740
rect 35950 6720 35970 6740
rect 35970 6720 36040 6740
rect 36040 6720 36070 6740
rect 35830 6700 36070 6720
rect 35830 6630 35860 6700
rect 35860 6630 35880 6700
rect 35880 6630 35950 6700
rect 35950 6630 35970 6700
rect 35970 6630 36040 6700
rect 36040 6630 36070 6700
rect 35830 6610 36070 6630
rect 35830 6540 35860 6610
rect 35860 6540 35880 6610
rect 35880 6540 35950 6610
rect 35950 6540 35970 6610
rect 35970 6540 36040 6610
rect 36040 6540 36070 6610
rect 35830 6520 36070 6540
rect 35830 6500 35860 6520
rect 35860 6500 35880 6520
rect 35880 6500 35950 6520
rect 35950 6500 35970 6520
rect 35970 6500 36040 6520
rect 36040 6500 36070 6520
rect 35830 6360 35860 6410
rect 35860 6360 35880 6410
rect 35880 6360 35950 6410
rect 35950 6360 35970 6410
rect 35970 6360 36040 6410
rect 36040 6360 36070 6410
rect 35830 6340 36070 6360
rect 35830 6270 35860 6340
rect 35860 6270 35880 6340
rect 35880 6270 35950 6340
rect 35950 6270 35970 6340
rect 35970 6270 36040 6340
rect 36040 6270 36070 6340
rect 35830 6250 36070 6270
rect 35830 6180 35860 6250
rect 35860 6180 35880 6250
rect 35880 6180 35950 6250
rect 35950 6180 35970 6250
rect 35970 6180 36040 6250
rect 36040 6180 36070 6250
rect 35830 6170 36070 6180
rect 35830 6070 36070 6080
rect 35830 6000 35860 6070
rect 35860 6000 35880 6070
rect 35880 6000 35950 6070
rect 35950 6000 35970 6070
rect 35970 6000 36040 6070
rect 36040 6000 36070 6070
rect 35830 5980 36070 6000
rect 35830 5910 35860 5980
rect 35860 5910 35880 5980
rect 35880 5910 35950 5980
rect 35950 5910 35970 5980
rect 35970 5910 36040 5980
rect 36040 5910 36070 5980
rect 35830 5890 36070 5910
rect 35830 5840 35860 5890
rect 35860 5840 35880 5890
rect 35880 5840 35950 5890
rect 35950 5840 35970 5890
rect 35970 5840 36040 5890
rect 36040 5840 36070 5890
rect 35830 5730 35860 5750
rect 35860 5730 35880 5750
rect 35880 5730 35950 5750
rect 35950 5730 35970 5750
rect 35970 5730 36040 5750
rect 36040 5730 36070 5750
rect 35830 5710 36070 5730
rect 35830 5640 35860 5710
rect 35860 5640 35880 5710
rect 35880 5640 35950 5710
rect 35950 5640 35970 5710
rect 35970 5640 36040 5710
rect 36040 5640 36070 5710
rect 35830 5620 36070 5640
rect 35830 5550 35860 5620
rect 35860 5550 35880 5620
rect 35880 5550 35950 5620
rect 35950 5550 35970 5620
rect 35970 5550 36040 5620
rect 36040 5550 36070 5620
rect 35830 5530 36070 5550
rect 35830 5510 35860 5530
rect 35860 5510 35880 5530
rect 35880 5510 35950 5530
rect 35950 5510 35970 5530
rect 35970 5510 36040 5530
rect 36040 5510 36070 5530
rect 35830 5370 35860 5420
rect 35860 5370 35880 5420
rect 35880 5370 35950 5420
rect 35950 5370 35970 5420
rect 35970 5370 36040 5420
rect 36040 5370 36070 5420
rect 35830 5350 36070 5370
rect 35830 5280 35860 5350
rect 35860 5280 35880 5350
rect 35880 5280 35950 5350
rect 35950 5280 35970 5350
rect 35970 5280 36040 5350
rect 36040 5280 36070 5350
rect 35830 5260 36070 5280
rect 35830 5190 35860 5260
rect 35860 5190 35880 5260
rect 35880 5190 35950 5260
rect 35950 5190 35970 5260
rect 35970 5190 36040 5260
rect 36040 5190 36070 5260
rect 35830 5180 36070 5190
rect 35830 5080 36070 5090
rect 35830 5010 35860 5080
rect 35860 5010 35880 5080
rect 35880 5010 35950 5080
rect 35950 5010 35970 5080
rect 35970 5010 36040 5080
rect 36040 5010 36070 5080
rect 35830 4990 36070 5010
rect 35830 4920 35860 4990
rect 35860 4920 35880 4990
rect 35880 4920 35950 4990
rect 35950 4920 35970 4990
rect 35970 4920 36040 4990
rect 36040 4920 36070 4990
rect 35830 4900 36070 4920
rect 35830 4850 35860 4900
rect 35860 4850 35880 4900
rect 35880 4850 35950 4900
rect 35950 4850 35970 4900
rect 35970 4850 36040 4900
rect 36040 4850 36070 4900
rect 35830 4740 35860 4760
rect 35860 4740 35880 4760
rect 35880 4740 35950 4760
rect 35950 4740 35970 4760
rect 35970 4740 36040 4760
rect 36040 4740 36070 4760
rect 35830 4720 36070 4740
rect 35830 4650 35860 4720
rect 35860 4650 35880 4720
rect 35880 4650 35950 4720
rect 35950 4650 35970 4720
rect 35970 4650 36040 4720
rect 36040 4650 36070 4720
rect 35830 4630 36070 4650
rect 35830 4560 35860 4630
rect 35860 4560 35880 4630
rect 35880 4560 35950 4630
rect 35950 4560 35970 4630
rect 35970 4560 36040 4630
rect 36040 4560 36070 4630
rect 35830 4540 36070 4560
rect 35830 4520 35860 4540
rect 35860 4520 35880 4540
rect 35880 4520 35950 4540
rect 35950 4520 35970 4540
rect 35970 4520 36040 4540
rect 36040 4520 36070 4540
rect 35830 4380 35860 4430
rect 35860 4380 35880 4430
rect 35880 4380 35950 4430
rect 35950 4380 35970 4430
rect 35970 4380 36040 4430
rect 36040 4380 36070 4430
rect 35830 4360 36070 4380
rect 35830 4290 35860 4360
rect 35860 4290 35880 4360
rect 35880 4290 35950 4360
rect 35950 4290 35970 4360
rect 35970 4290 36040 4360
rect 36040 4290 36070 4360
rect 35830 4270 36070 4290
rect 35830 4200 35860 4270
rect 35860 4200 35880 4270
rect 35880 4200 35950 4270
rect 35950 4200 35970 4270
rect 35970 4200 36040 4270
rect 36040 4200 36070 4270
rect 35830 4190 36070 4200
rect 35830 4050 36070 4060
rect 35830 3980 35860 4050
rect 35860 3980 35880 4050
rect 35880 3980 35950 4050
rect 35950 3980 35970 4050
rect 35970 3980 36040 4050
rect 36040 3980 36070 4050
rect 35830 3960 36070 3980
rect 35830 3890 35860 3960
rect 35860 3890 35880 3960
rect 35880 3890 35950 3960
rect 35950 3890 35970 3960
rect 35970 3890 36040 3960
rect 36040 3890 36070 3960
rect 35830 3870 36070 3890
rect 35830 3820 35860 3870
rect 35860 3820 35880 3870
rect 35880 3820 35950 3870
rect 35950 3820 35970 3870
rect 35970 3820 36040 3870
rect 36040 3820 36070 3870
rect 35830 3710 35860 3730
rect 35860 3710 35880 3730
rect 35880 3710 35950 3730
rect 35950 3710 35970 3730
rect 35970 3710 36040 3730
rect 36040 3710 36070 3730
rect 35830 3690 36070 3710
rect 35830 3620 35860 3690
rect 35860 3620 35880 3690
rect 35880 3620 35950 3690
rect 35950 3620 35970 3690
rect 35970 3620 36040 3690
rect 36040 3620 36070 3690
rect 35830 3600 36070 3620
rect 35830 3530 35860 3600
rect 35860 3530 35880 3600
rect 35880 3530 35950 3600
rect 35950 3530 35970 3600
rect 35970 3530 36040 3600
rect 36040 3530 36070 3600
rect 35830 3510 36070 3530
rect 35830 3490 35860 3510
rect 35860 3490 35880 3510
rect 35880 3490 35950 3510
rect 35950 3490 35970 3510
rect 35970 3490 36040 3510
rect 36040 3490 36070 3510
rect 35830 3350 35860 3400
rect 35860 3350 35880 3400
rect 35880 3350 35950 3400
rect 35950 3350 35970 3400
rect 35970 3350 36040 3400
rect 36040 3350 36070 3400
rect 35830 3330 36070 3350
rect 35830 3260 35860 3330
rect 35860 3260 35880 3330
rect 35880 3260 35950 3330
rect 35950 3260 35970 3330
rect 35970 3260 36040 3330
rect 36040 3260 36070 3330
rect 35830 3240 36070 3260
rect 35830 3170 35860 3240
rect 35860 3170 35880 3240
rect 35880 3170 35950 3240
rect 35950 3170 35970 3240
rect 35970 3170 36040 3240
rect 36040 3170 36070 3240
rect 35830 3160 36070 3170
rect 35830 3060 36070 3070
rect 35830 2990 35860 3060
rect 35860 2990 35880 3060
rect 35880 2990 35950 3060
rect 35950 2990 35970 3060
rect 35970 2990 36040 3060
rect 36040 2990 36070 3060
rect 35830 2970 36070 2990
rect 35830 2900 35860 2970
rect 35860 2900 35880 2970
rect 35880 2900 35950 2970
rect 35950 2900 35970 2970
rect 35970 2900 36040 2970
rect 36040 2900 36070 2970
rect 35830 2880 36070 2900
rect 35830 2830 35860 2880
rect 35860 2830 35880 2880
rect 35880 2830 35950 2880
rect 35950 2830 35970 2880
rect 35970 2830 36040 2880
rect 36040 2830 36070 2880
rect 35830 2720 35860 2740
rect 35860 2720 35880 2740
rect 35880 2720 35950 2740
rect 35950 2720 35970 2740
rect 35970 2720 36040 2740
rect 36040 2720 36070 2740
rect 35830 2700 36070 2720
rect 35830 2630 35860 2700
rect 35860 2630 35880 2700
rect 35880 2630 35950 2700
rect 35950 2630 35970 2700
rect 35970 2630 36040 2700
rect 36040 2630 36070 2700
rect 35830 2610 36070 2630
rect 35830 2540 35860 2610
rect 35860 2540 35880 2610
rect 35880 2540 35950 2610
rect 35950 2540 35970 2610
rect 35970 2540 36040 2610
rect 36040 2540 36070 2610
rect 35830 2520 36070 2540
rect 35830 2500 35860 2520
rect 35860 2500 35880 2520
rect 35880 2500 35950 2520
rect 35950 2500 35970 2520
rect 35970 2500 36040 2520
rect 36040 2500 36070 2520
rect 35830 2360 35860 2410
rect 35860 2360 35880 2410
rect 35880 2360 35950 2410
rect 35950 2360 35970 2410
rect 35970 2360 36040 2410
rect 36040 2360 36070 2410
rect 35830 2340 36070 2360
rect 35830 2270 35860 2340
rect 35860 2270 35880 2340
rect 35880 2270 35950 2340
rect 35950 2270 35970 2340
rect 35970 2270 36040 2340
rect 36040 2270 36070 2340
rect 35830 2250 36070 2270
rect 35830 2180 35860 2250
rect 35860 2180 35880 2250
rect 35880 2180 35950 2250
rect 35950 2180 35970 2250
rect 35970 2180 36040 2250
rect 36040 2180 36070 2250
rect 35830 2170 36070 2180
rect 35830 2070 36070 2080
rect 35830 2000 35860 2070
rect 35860 2000 35880 2070
rect 35880 2000 35950 2070
rect 35950 2000 35970 2070
rect 35970 2000 36040 2070
rect 36040 2000 36070 2070
rect 35830 1980 36070 2000
rect 35830 1910 35860 1980
rect 35860 1910 35880 1980
rect 35880 1910 35950 1980
rect 35950 1910 35970 1980
rect 35970 1910 36040 1980
rect 36040 1910 36070 1980
rect 35830 1890 36070 1910
rect 35830 1840 35860 1890
rect 35860 1840 35880 1890
rect 35880 1840 35950 1890
rect 35950 1840 35970 1890
rect 35970 1840 36040 1890
rect 36040 1840 36070 1890
rect 35830 1730 35860 1750
rect 35860 1730 35880 1750
rect 35880 1730 35950 1750
rect 35950 1730 35970 1750
rect 35970 1730 36040 1750
rect 36040 1730 36070 1750
rect 35830 1710 36070 1730
rect 35830 1640 35860 1710
rect 35860 1640 35880 1710
rect 35880 1640 35950 1710
rect 35950 1640 35970 1710
rect 35970 1640 36040 1710
rect 36040 1640 36070 1710
rect 35830 1620 36070 1640
rect 35830 1550 35860 1620
rect 35860 1550 35880 1620
rect 35880 1550 35950 1620
rect 35950 1550 35970 1620
rect 35970 1550 36040 1620
rect 36040 1550 36070 1620
rect 35830 1530 36070 1550
rect 35830 1510 35860 1530
rect 35860 1510 35880 1530
rect 35880 1510 35950 1530
rect 35950 1510 35970 1530
rect 35970 1510 36040 1530
rect 36040 1510 36070 1530
rect 35830 1370 35860 1420
rect 35860 1370 35880 1420
rect 35880 1370 35950 1420
rect 35950 1370 35970 1420
rect 35970 1370 36040 1420
rect 36040 1370 36070 1420
rect 35830 1350 36070 1370
rect 35830 1280 35860 1350
rect 35860 1280 35880 1350
rect 35880 1280 35950 1350
rect 35950 1280 35970 1350
rect 35970 1280 36040 1350
rect 36040 1280 36070 1350
rect 35830 1260 36070 1280
rect 35830 1190 35860 1260
rect 35860 1190 35880 1260
rect 35880 1190 35950 1260
rect 35950 1190 35970 1260
rect 35970 1190 36040 1260
rect 36040 1190 36070 1260
rect 35830 1180 36070 1190
rect 20080 -3760 20140 -3690
rect 20140 -3760 20180 -3690
rect 20180 -3760 20250 -3690
rect 20250 -3760 20290 -3690
rect 20290 -3760 20360 -3690
rect 20360 -3760 20400 -3690
rect 20400 -3760 20450 -3690
rect 20080 -3800 20450 -3760
rect 20080 -3870 20140 -3800
rect 20140 -3870 20180 -3800
rect 20180 -3870 20250 -3800
rect 20250 -3870 20290 -3800
rect 20290 -3870 20360 -3800
rect 20360 -3870 20400 -3800
rect 20400 -3870 20450 -3800
rect 20080 -3930 20450 -3870
rect 24560 -3760 24620 -3690
rect 24620 -3760 24660 -3690
rect 24660 -3760 24730 -3690
rect 24730 -3760 24770 -3690
rect 24770 -3760 24840 -3690
rect 24840 -3760 24880 -3690
rect 24880 -3760 24930 -3690
rect 24560 -3800 24930 -3760
rect 24560 -3870 24620 -3800
rect 24620 -3870 24660 -3800
rect 24660 -3870 24730 -3800
rect 24730 -3870 24770 -3800
rect 24770 -3870 24840 -3800
rect 24840 -3870 24880 -3800
rect 24880 -3870 24930 -3800
rect 24560 -3930 24930 -3870
rect -120 -7700 -90 -7650
rect -90 -7700 -70 -7650
rect -70 -7700 0 -7650
rect 0 -7700 20 -7650
rect 20 -7700 90 -7650
rect 90 -7700 120 -7650
rect -120 -7720 120 -7700
rect -120 -7790 -90 -7720
rect -90 -7790 -70 -7720
rect -70 -7790 0 -7720
rect 0 -7790 20 -7720
rect 20 -7790 90 -7720
rect 90 -7790 120 -7720
rect -120 -7810 120 -7790
rect -120 -7880 -90 -7810
rect -90 -7880 -70 -7810
rect -70 -7880 0 -7810
rect 0 -7880 20 -7810
rect 20 -7880 90 -7810
rect 90 -7880 120 -7810
rect -120 -7890 120 -7880
rect -120 -7990 120 -7980
rect -120 -8060 -90 -7990
rect -90 -8060 -70 -7990
rect -70 -8060 0 -7990
rect 0 -8060 20 -7990
rect 20 -8060 90 -7990
rect 90 -8060 120 -7990
rect -120 -8080 120 -8060
rect -120 -8150 -90 -8080
rect -90 -8150 -70 -8080
rect -70 -8150 0 -8080
rect 0 -8150 20 -8080
rect 20 -8150 90 -8080
rect 90 -8150 120 -8080
rect -120 -8170 120 -8150
rect -120 -8220 -90 -8170
rect -90 -8220 -70 -8170
rect -70 -8220 0 -8170
rect 0 -8220 20 -8170
rect 20 -8220 90 -8170
rect 90 -8220 120 -8170
rect -120 -8330 -90 -8310
rect -90 -8330 -70 -8310
rect -70 -8330 0 -8310
rect 0 -8330 20 -8310
rect 20 -8330 90 -8310
rect 90 -8330 120 -8310
rect -120 -8350 120 -8330
rect -120 -8420 -90 -8350
rect -90 -8420 -70 -8350
rect -70 -8420 0 -8350
rect 0 -8420 20 -8350
rect 20 -8420 90 -8350
rect 90 -8420 120 -8350
rect -120 -8440 120 -8420
rect -120 -8510 -90 -8440
rect -90 -8510 -70 -8440
rect -70 -8510 0 -8440
rect 0 -8510 20 -8440
rect 20 -8510 90 -8440
rect 90 -8510 120 -8440
rect -120 -8530 120 -8510
rect -120 -8550 -90 -8530
rect -90 -8550 -70 -8530
rect -70 -8550 0 -8530
rect 0 -8550 20 -8530
rect 20 -8550 90 -8530
rect 90 -8550 120 -8530
rect -120 -8690 -90 -8640
rect -90 -8690 -70 -8640
rect -70 -8690 0 -8640
rect 0 -8690 20 -8640
rect 20 -8690 90 -8640
rect 90 -8690 120 -8640
rect -120 -8710 120 -8690
rect -120 -8780 -90 -8710
rect -90 -8780 -70 -8710
rect -70 -8780 0 -8710
rect 0 -8780 20 -8710
rect 20 -8780 90 -8710
rect 90 -8780 120 -8710
rect -120 -8800 120 -8780
rect -120 -8870 -90 -8800
rect -90 -8870 -70 -8800
rect -70 -8870 0 -8800
rect 0 -8870 20 -8800
rect 20 -8870 90 -8800
rect 90 -8870 120 -8800
rect -120 -8880 120 -8870
rect 19250 -8630 19300 -8570
rect 19300 -8630 19330 -8570
rect 19330 -8630 19400 -8570
rect 19400 -8630 19430 -8570
rect 19430 -8630 19490 -8570
rect 19250 -8660 19490 -8630
rect 19250 -8730 19300 -8660
rect 19300 -8730 19330 -8660
rect 19330 -8730 19400 -8660
rect 19400 -8730 19430 -8660
rect 19430 -8730 19490 -8660
rect 19250 -8760 19490 -8730
rect 19250 -8810 19300 -8760
rect 19300 -8810 19330 -8760
rect 19330 -8810 19400 -8760
rect 19400 -8810 19430 -8760
rect 19430 -8810 19490 -8760
rect 1260 -10410 1330 -10340
rect 1330 -10410 1370 -10340
rect 1370 -10410 1440 -10340
rect 1440 -10410 1480 -10340
rect 1480 -10410 1500 -10340
rect 1590 -10410 1660 -10340
rect 1660 -10410 1700 -10340
rect 1700 -10410 1770 -10340
rect 1770 -10410 1810 -10340
rect 1810 -10410 1830 -10340
rect 1930 -10410 1990 -10340
rect 1990 -10410 2030 -10340
rect 2030 -10410 2100 -10340
rect 2100 -10410 2140 -10340
rect 2140 -10410 2170 -10340
rect 2260 -10410 2320 -10340
rect 2320 -10410 2360 -10340
rect 2360 -10410 2430 -10340
rect 2430 -10410 2470 -10340
rect 2470 -10410 2500 -10340
rect 1260 -10450 1500 -10410
rect 1590 -10450 1830 -10410
rect 1930 -10450 2170 -10410
rect 2260 -10450 2500 -10410
rect 1260 -10520 1330 -10450
rect 1330 -10520 1370 -10450
rect 1370 -10520 1440 -10450
rect 1440 -10520 1480 -10450
rect 1480 -10520 1500 -10450
rect 1590 -10520 1660 -10450
rect 1660 -10520 1700 -10450
rect 1700 -10520 1770 -10450
rect 1770 -10520 1810 -10450
rect 1810 -10520 1830 -10450
rect 1930 -10520 1990 -10450
rect 1990 -10520 2030 -10450
rect 2030 -10520 2100 -10450
rect 2100 -10520 2140 -10450
rect 2140 -10520 2170 -10450
rect 2260 -10520 2320 -10450
rect 2320 -10520 2360 -10450
rect 2360 -10520 2430 -10450
rect 2430 -10520 2470 -10450
rect 2470 -10520 2500 -10450
rect 1260 -10580 1500 -10520
rect 1590 -10580 1830 -10520
rect 1930 -10580 2170 -10520
rect 2260 -10580 2500 -10520
rect 12400 -10440 12470 -10370
rect 12470 -10440 12510 -10370
rect 12510 -10440 12580 -10370
rect 12580 -10440 12620 -10370
rect 12620 -10440 12640 -10370
rect 12730 -10440 12800 -10370
rect 12800 -10440 12840 -10370
rect 12840 -10440 12910 -10370
rect 12910 -10440 12950 -10370
rect 12950 -10440 12970 -10370
rect 13070 -10440 13130 -10370
rect 13130 -10440 13170 -10370
rect 13170 -10440 13240 -10370
rect 13240 -10440 13280 -10370
rect 13280 -10440 13310 -10370
rect 13400 -10440 13460 -10370
rect 13460 -10440 13500 -10370
rect 13500 -10440 13570 -10370
rect 13570 -10440 13610 -10370
rect 13610 -10440 13640 -10370
rect 12400 -10480 12640 -10440
rect 12730 -10480 12970 -10440
rect 13070 -10480 13310 -10440
rect 13400 -10480 13640 -10440
rect 12400 -10550 12470 -10480
rect 12470 -10550 12510 -10480
rect 12510 -10550 12580 -10480
rect 12580 -10550 12620 -10480
rect 12620 -10550 12640 -10480
rect 12730 -10550 12800 -10480
rect 12800 -10550 12840 -10480
rect 12840 -10550 12910 -10480
rect 12910 -10550 12950 -10480
rect 12950 -10550 12970 -10480
rect 13070 -10550 13130 -10480
rect 13130 -10550 13170 -10480
rect 13170 -10550 13240 -10480
rect 13240 -10550 13280 -10480
rect 13280 -10550 13310 -10480
rect 13400 -10550 13460 -10480
rect 13460 -10550 13500 -10480
rect 13500 -10550 13570 -10480
rect 13570 -10550 13610 -10480
rect 13610 -10550 13640 -10480
rect 12400 -10610 12640 -10550
rect 12730 -10610 12970 -10550
rect 13070 -10610 13310 -10550
rect 13400 -10610 13640 -10550
rect 35830 150 35860 170
rect 35860 150 35880 170
rect 35880 150 35950 170
rect 35950 150 35970 170
rect 35970 150 36040 170
rect 36040 150 36070 170
rect 35830 130 36070 150
rect 35830 60 35860 130
rect 35860 60 35880 130
rect 35880 60 35950 130
rect 35950 60 35970 130
rect 35970 60 36040 130
rect 36040 60 36070 130
rect 35830 40 36070 60
rect 35830 -30 35860 40
rect 35860 -30 35880 40
rect 35880 -30 35950 40
rect 35950 -30 35970 40
rect 35970 -30 36040 40
rect 36040 -30 36070 40
rect 35830 -50 36070 -30
rect 35830 -70 35860 -50
rect 35860 -70 35880 -50
rect 35880 -70 35950 -50
rect 35950 -70 35970 -50
rect 35970 -70 36040 -50
rect 36040 -70 36070 -50
rect 35830 -210 35860 -160
rect 35860 -210 35880 -160
rect 35880 -210 35950 -160
rect 35950 -210 35970 -160
rect 35970 -210 36040 -160
rect 36040 -210 36070 -160
rect 35830 -230 36070 -210
rect 35830 -300 35860 -230
rect 35860 -300 35880 -230
rect 35880 -300 35950 -230
rect 35950 -300 35970 -230
rect 35970 -300 36040 -230
rect 36040 -300 36070 -230
rect 35830 -320 36070 -300
rect 35830 -390 35860 -320
rect 35860 -390 35880 -320
rect 35880 -390 35950 -320
rect 35950 -390 35970 -320
rect 35970 -390 36040 -320
rect 36040 -390 36070 -320
rect 35830 -400 36070 -390
rect 35830 -540 36070 -530
rect 35830 -610 35860 -540
rect 35860 -610 35880 -540
rect 35880 -610 35950 -540
rect 35950 -610 35970 -540
rect 35970 -610 36040 -540
rect 36040 -610 36070 -540
rect 35830 -630 36070 -610
rect 35830 -700 35860 -630
rect 35860 -700 35880 -630
rect 35880 -700 35950 -630
rect 35950 -700 35970 -630
rect 35970 -700 36040 -630
rect 36040 -700 36070 -630
rect 35830 -720 36070 -700
rect 35830 -770 35860 -720
rect 35860 -770 35880 -720
rect 35880 -770 35950 -720
rect 35950 -770 35970 -720
rect 35970 -770 36040 -720
rect 36040 -770 36070 -720
rect 35830 -880 35860 -860
rect 35860 -880 35880 -860
rect 35880 -880 35950 -860
rect 35950 -880 35970 -860
rect 35970 -880 36040 -860
rect 36040 -880 36070 -860
rect 35830 -900 36070 -880
rect 35830 -970 35860 -900
rect 35860 -970 35880 -900
rect 35880 -970 35950 -900
rect 35950 -970 35970 -900
rect 35970 -970 36040 -900
rect 36040 -970 36070 -900
rect 35830 -990 36070 -970
rect 35830 -1060 35860 -990
rect 35860 -1060 35880 -990
rect 35880 -1060 35950 -990
rect 35950 -1060 35970 -990
rect 35970 -1060 36040 -990
rect 36040 -1060 36070 -990
rect 35830 -1080 36070 -1060
rect 35830 -1100 35860 -1080
rect 35860 -1100 35880 -1080
rect 35880 -1100 35950 -1080
rect 35950 -1100 35970 -1080
rect 35970 -1100 36040 -1080
rect 36040 -1100 36070 -1080
rect 35830 -1240 35860 -1190
rect 35860 -1240 35880 -1190
rect 35880 -1240 35950 -1190
rect 35950 -1240 35970 -1190
rect 35970 -1240 36040 -1190
rect 36040 -1240 36070 -1190
rect 35830 -1260 36070 -1240
rect 35830 -1330 35860 -1260
rect 35860 -1330 35880 -1260
rect 35880 -1330 35950 -1260
rect 35950 -1330 35970 -1260
rect 35970 -1330 36040 -1260
rect 36040 -1330 36070 -1260
rect 35830 -1350 36070 -1330
rect 35830 -1420 35860 -1350
rect 35860 -1420 35880 -1350
rect 35880 -1420 35950 -1350
rect 35950 -1420 35970 -1350
rect 35970 -1420 36040 -1350
rect 36040 -1420 36070 -1350
rect 35830 -1430 36070 -1420
rect 35830 -1530 36070 -1520
rect 35830 -1600 35860 -1530
rect 35860 -1600 35880 -1530
rect 35880 -1600 35950 -1530
rect 35950 -1600 35970 -1530
rect 35970 -1600 36040 -1530
rect 36040 -1600 36070 -1530
rect 35830 -1620 36070 -1600
rect 35830 -1690 35860 -1620
rect 35860 -1690 35880 -1620
rect 35880 -1690 35950 -1620
rect 35950 -1690 35970 -1620
rect 35970 -1690 36040 -1620
rect 36040 -1690 36070 -1620
rect 35830 -1710 36070 -1690
rect 35830 -1760 35860 -1710
rect 35860 -1760 35880 -1710
rect 35880 -1760 35950 -1710
rect 35950 -1760 35970 -1710
rect 35970 -1760 36040 -1710
rect 36040 -1760 36070 -1710
rect 35830 -1870 35860 -1850
rect 35860 -1870 35880 -1850
rect 35880 -1870 35950 -1850
rect 35950 -1870 35970 -1850
rect 35970 -1870 36040 -1850
rect 36040 -1870 36070 -1850
rect 35830 -1890 36070 -1870
rect 35830 -1960 35860 -1890
rect 35860 -1960 35880 -1890
rect 35880 -1960 35950 -1890
rect 35950 -1960 35970 -1890
rect 35970 -1960 36040 -1890
rect 36040 -1960 36070 -1890
rect 35830 -1980 36070 -1960
rect 35830 -2050 35860 -1980
rect 35860 -2050 35880 -1980
rect 35880 -2050 35950 -1980
rect 35950 -2050 35970 -1980
rect 35970 -2050 36040 -1980
rect 36040 -2050 36070 -1980
rect 35830 -2070 36070 -2050
rect 35830 -2090 35860 -2070
rect 35860 -2090 35880 -2070
rect 35880 -2090 35950 -2070
rect 35950 -2090 35970 -2070
rect 35970 -2090 36040 -2070
rect 36040 -2090 36070 -2070
rect 35830 -2230 35860 -2180
rect 35860 -2230 35880 -2180
rect 35880 -2230 35950 -2180
rect 35950 -2230 35970 -2180
rect 35970 -2230 36040 -2180
rect 36040 -2230 36070 -2180
rect 35830 -2250 36070 -2230
rect 35830 -2320 35860 -2250
rect 35860 -2320 35880 -2250
rect 35880 -2320 35950 -2250
rect 35950 -2320 35970 -2250
rect 35970 -2320 36040 -2250
rect 36040 -2320 36070 -2250
rect 35830 -2340 36070 -2320
rect 35830 -2410 35860 -2340
rect 35860 -2410 35880 -2340
rect 35880 -2410 35950 -2340
rect 35950 -2410 35970 -2340
rect 35970 -2410 36040 -2340
rect 36040 -2410 36070 -2340
rect 35830 -2420 36070 -2410
rect 35830 -2520 36070 -2510
rect 35830 -2590 35860 -2520
rect 35860 -2590 35880 -2520
rect 35880 -2590 35950 -2520
rect 35950 -2590 35970 -2520
rect 35970 -2590 36040 -2520
rect 36040 -2590 36070 -2520
rect 35830 -2610 36070 -2590
rect 35830 -2680 35860 -2610
rect 35860 -2680 35880 -2610
rect 35880 -2680 35950 -2610
rect 35950 -2680 35970 -2610
rect 35970 -2680 36040 -2610
rect 36040 -2680 36070 -2610
rect 35830 -2700 36070 -2680
rect 35830 -2750 35860 -2700
rect 35860 -2750 35880 -2700
rect 35880 -2750 35950 -2700
rect 35950 -2750 35970 -2700
rect 35970 -2750 36040 -2700
rect 36040 -2750 36070 -2700
rect 35830 -2860 35860 -2840
rect 35860 -2860 35880 -2840
rect 35880 -2860 35950 -2840
rect 35950 -2860 35970 -2840
rect 35970 -2860 36040 -2840
rect 36040 -2860 36070 -2840
rect 35830 -2880 36070 -2860
rect 35830 -2950 35860 -2880
rect 35860 -2950 35880 -2880
rect 35880 -2950 35950 -2880
rect 35950 -2950 35970 -2880
rect 35970 -2950 36040 -2880
rect 36040 -2950 36070 -2880
rect 35830 -2970 36070 -2950
rect 35830 -3040 35860 -2970
rect 35860 -3040 35880 -2970
rect 35880 -3040 35950 -2970
rect 35950 -3040 35970 -2970
rect 35970 -3040 36040 -2970
rect 36040 -3040 36070 -2970
rect 35830 -3060 36070 -3040
rect 35830 -3080 35860 -3060
rect 35860 -3080 35880 -3060
rect 35880 -3080 35950 -3060
rect 35950 -3080 35970 -3060
rect 35970 -3080 36040 -3060
rect 36040 -3080 36070 -3060
rect 35830 -3220 35860 -3170
rect 35860 -3220 35880 -3170
rect 35880 -3220 35950 -3170
rect 35950 -3220 35970 -3170
rect 35970 -3220 36040 -3170
rect 36040 -3220 36070 -3170
rect 35830 -3240 36070 -3220
rect 35830 -3310 35860 -3240
rect 35860 -3310 35880 -3240
rect 35880 -3310 35950 -3240
rect 35950 -3310 35970 -3240
rect 35970 -3310 36040 -3240
rect 36040 -3310 36070 -3240
rect 35830 -3330 36070 -3310
rect 35830 -3400 35860 -3330
rect 35860 -3400 35880 -3330
rect 35880 -3400 35950 -3330
rect 35950 -3400 35970 -3330
rect 35970 -3400 36040 -3330
rect 36040 -3400 36070 -3330
rect 35830 -3410 36070 -3400
rect 35830 -3550 36070 -3540
rect 35830 -3620 35860 -3550
rect 35860 -3620 35880 -3550
rect 35880 -3620 35950 -3550
rect 35950 -3620 35970 -3550
rect 35970 -3620 36040 -3550
rect 36040 -3620 36070 -3550
rect 35830 -3640 36070 -3620
rect 35830 -3710 35860 -3640
rect 35860 -3710 35880 -3640
rect 35880 -3710 35950 -3640
rect 35950 -3710 35970 -3640
rect 35970 -3710 36040 -3640
rect 36040 -3710 36070 -3640
rect 35830 -3730 36070 -3710
rect 35830 -3780 35860 -3730
rect 35860 -3780 35880 -3730
rect 35880 -3780 35950 -3730
rect 35950 -3780 35970 -3730
rect 35970 -3780 36040 -3730
rect 36040 -3780 36070 -3730
rect 35830 -3890 35860 -3870
rect 35860 -3890 35880 -3870
rect 35880 -3890 35950 -3870
rect 35950 -3890 35970 -3870
rect 35970 -3890 36040 -3870
rect 36040 -3890 36070 -3870
rect 35830 -3910 36070 -3890
rect 35830 -3980 35860 -3910
rect 35860 -3980 35880 -3910
rect 35880 -3980 35950 -3910
rect 35950 -3980 35970 -3910
rect 35970 -3980 36040 -3910
rect 36040 -3980 36070 -3910
rect 35830 -4000 36070 -3980
rect 35830 -4070 35860 -4000
rect 35860 -4070 35880 -4000
rect 35880 -4070 35950 -4000
rect 35950 -4070 35970 -4000
rect 35970 -4070 36040 -4000
rect 36040 -4070 36070 -4000
rect 35830 -4090 36070 -4070
rect 35830 -4110 35860 -4090
rect 35860 -4110 35880 -4090
rect 35880 -4110 35950 -4090
rect 35950 -4110 35970 -4090
rect 35970 -4110 36040 -4090
rect 36040 -4110 36070 -4090
rect 35830 -4250 35860 -4200
rect 35860 -4250 35880 -4200
rect 35880 -4250 35950 -4200
rect 35950 -4250 35970 -4200
rect 35970 -4250 36040 -4200
rect 36040 -4250 36070 -4200
rect 35830 -4270 36070 -4250
rect 35830 -4340 35860 -4270
rect 35860 -4340 35880 -4270
rect 35880 -4340 35950 -4270
rect 35950 -4340 35970 -4270
rect 35970 -4340 36040 -4270
rect 36040 -4340 36070 -4270
rect 35830 -4360 36070 -4340
rect 35830 -4430 35860 -4360
rect 35860 -4430 35880 -4360
rect 35880 -4430 35950 -4360
rect 35950 -4430 35970 -4360
rect 35970 -4430 36040 -4360
rect 36040 -4430 36070 -4360
rect 35830 -4440 36070 -4430
rect 35830 -4540 36070 -4530
rect 35830 -4610 35860 -4540
rect 35860 -4610 35880 -4540
rect 35880 -4610 35950 -4540
rect 35950 -4610 35970 -4540
rect 35970 -4610 36040 -4540
rect 36040 -4610 36070 -4540
rect 35830 -4630 36070 -4610
rect 35830 -4700 35860 -4630
rect 35860 -4700 35880 -4630
rect 35880 -4700 35950 -4630
rect 35950 -4700 35970 -4630
rect 35970 -4700 36040 -4630
rect 36040 -4700 36070 -4630
rect 35830 -4720 36070 -4700
rect 35830 -4770 35860 -4720
rect 35860 -4770 35880 -4720
rect 35880 -4770 35950 -4720
rect 35950 -4770 35970 -4720
rect 35970 -4770 36040 -4720
rect 36040 -4770 36070 -4720
rect 35830 -4880 35860 -4860
rect 35860 -4880 35880 -4860
rect 35880 -4880 35950 -4860
rect 35950 -4880 35970 -4860
rect 35970 -4880 36040 -4860
rect 36040 -4880 36070 -4860
rect 35830 -4900 36070 -4880
rect 35830 -4970 35860 -4900
rect 35860 -4970 35880 -4900
rect 35880 -4970 35950 -4900
rect 35950 -4970 35970 -4900
rect 35970 -4970 36040 -4900
rect 36040 -4970 36070 -4900
rect 35830 -4990 36070 -4970
rect 35830 -5060 35860 -4990
rect 35860 -5060 35880 -4990
rect 35880 -5060 35950 -4990
rect 35950 -5060 35970 -4990
rect 35970 -5060 36040 -4990
rect 36040 -5060 36070 -4990
rect 35830 -5080 36070 -5060
rect 35830 -5100 35860 -5080
rect 35860 -5100 35880 -5080
rect 35880 -5100 35950 -5080
rect 35950 -5100 35970 -5080
rect 35970 -5100 36040 -5080
rect 36040 -5100 36070 -5080
rect 35830 -5240 35860 -5190
rect 35860 -5240 35880 -5190
rect 35880 -5240 35950 -5190
rect 35950 -5240 35970 -5190
rect 35970 -5240 36040 -5190
rect 36040 -5240 36070 -5190
rect 35830 -5260 36070 -5240
rect 35830 -5330 35860 -5260
rect 35860 -5330 35880 -5260
rect 35880 -5330 35950 -5260
rect 35950 -5330 35970 -5260
rect 35970 -5330 36040 -5260
rect 36040 -5330 36070 -5260
rect 35830 -5350 36070 -5330
rect 35830 -5420 35860 -5350
rect 35860 -5420 35880 -5350
rect 35880 -5420 35950 -5350
rect 35950 -5420 35970 -5350
rect 35970 -5420 36040 -5350
rect 36040 -5420 36070 -5350
rect 35830 -5430 36070 -5420
rect 35830 -5530 36070 -5520
rect 35830 -5600 35860 -5530
rect 35860 -5600 35880 -5530
rect 35880 -5600 35950 -5530
rect 35950 -5600 35970 -5530
rect 35970 -5600 36040 -5530
rect 36040 -5600 36070 -5530
rect 35830 -5620 36070 -5600
rect 35830 -5690 35860 -5620
rect 35860 -5690 35880 -5620
rect 35880 -5690 35950 -5620
rect 35950 -5690 35970 -5620
rect 35970 -5690 36040 -5620
rect 36040 -5690 36070 -5620
rect 35830 -5710 36070 -5690
rect 35830 -5760 35860 -5710
rect 35860 -5760 35880 -5710
rect 35880 -5760 35950 -5710
rect 35950 -5760 35970 -5710
rect 35970 -5760 36040 -5710
rect 36040 -5760 36070 -5710
rect 35830 -5870 35860 -5850
rect 35860 -5870 35880 -5850
rect 35880 -5870 35950 -5850
rect 35950 -5870 35970 -5850
rect 35970 -5870 36040 -5850
rect 36040 -5870 36070 -5850
rect 35830 -5890 36070 -5870
rect 35830 -5960 35860 -5890
rect 35860 -5960 35880 -5890
rect 35880 -5960 35950 -5890
rect 35950 -5960 35970 -5890
rect 35970 -5960 36040 -5890
rect 36040 -5960 36070 -5890
rect 35830 -5980 36070 -5960
rect 35830 -6050 35860 -5980
rect 35860 -6050 35880 -5980
rect 35880 -6050 35950 -5980
rect 35950 -6050 35970 -5980
rect 35970 -6050 36040 -5980
rect 36040 -6050 36070 -5980
rect 35830 -6070 36070 -6050
rect 35830 -6090 35860 -6070
rect 35860 -6090 35880 -6070
rect 35880 -6090 35950 -6070
rect 35950 -6090 35970 -6070
rect 35970 -6090 36040 -6070
rect 36040 -6090 36070 -6070
rect 35830 -6230 35860 -6180
rect 35860 -6230 35880 -6180
rect 35880 -6230 35950 -6180
rect 35950 -6230 35970 -6180
rect 35970 -6230 36040 -6180
rect 36040 -6230 36070 -6180
rect 35830 -6250 36070 -6230
rect 35830 -6320 35860 -6250
rect 35860 -6320 35880 -6250
rect 35880 -6320 35950 -6250
rect 35950 -6320 35970 -6250
rect 35970 -6320 36040 -6250
rect 36040 -6320 36070 -6250
rect 35830 -6340 36070 -6320
rect 35830 -6410 35860 -6340
rect 35860 -6410 35880 -6340
rect 35880 -6410 35950 -6340
rect 35950 -6410 35970 -6340
rect 35970 -6410 36040 -6340
rect 36040 -6410 36070 -6340
rect 35830 -6420 36070 -6410
rect 2390 -12300 2630 -12240
rect 2720 -12300 2960 -12240
rect 3060 -12300 3300 -12240
rect 3390 -12300 3630 -12240
rect 2390 -12370 2420 -12300
rect 2420 -12370 2460 -12300
rect 2460 -12370 2530 -12300
rect 2530 -12370 2570 -12300
rect 2570 -12370 2630 -12300
rect 2720 -12370 2750 -12300
rect 2750 -12370 2790 -12300
rect 2790 -12370 2860 -12300
rect 2860 -12370 2900 -12300
rect 2900 -12370 2960 -12300
rect 3060 -12370 3080 -12300
rect 3080 -12370 3120 -12300
rect 3120 -12370 3190 -12300
rect 3190 -12370 3230 -12300
rect 3230 -12370 3300 -12300
rect 3390 -12370 3410 -12300
rect 3410 -12370 3450 -12300
rect 3450 -12370 3520 -12300
rect 3520 -12370 3560 -12300
rect 3560 -12370 3630 -12300
rect 2390 -12410 2630 -12370
rect 2720 -12410 2960 -12370
rect 3060 -12410 3300 -12370
rect 3390 -12410 3630 -12370
rect 2390 -12480 2420 -12410
rect 2420 -12480 2460 -12410
rect 2460 -12480 2530 -12410
rect 2530 -12480 2570 -12410
rect 2570 -12480 2630 -12410
rect 2720 -12480 2750 -12410
rect 2750 -12480 2790 -12410
rect 2790 -12480 2860 -12410
rect 2860 -12480 2900 -12410
rect 2900 -12480 2960 -12410
rect 3060 -12480 3080 -12410
rect 3080 -12480 3120 -12410
rect 3120 -12480 3190 -12410
rect 3190 -12480 3230 -12410
rect 3230 -12480 3300 -12410
rect 3390 -12480 3410 -12410
rect 3410 -12480 3450 -12410
rect 3450 -12480 3520 -12410
rect 3520 -12480 3560 -12410
rect 3560 -12480 3630 -12410
rect 11270 -12300 11510 -12240
rect 11600 -12300 11840 -12240
rect 11940 -12300 12180 -12240
rect 12270 -12300 12510 -12240
rect 11270 -12370 11300 -12300
rect 11300 -12370 11340 -12300
rect 11340 -12370 11410 -12300
rect 11410 -12370 11450 -12300
rect 11450 -12370 11510 -12300
rect 11600 -12370 11630 -12300
rect 11630 -12370 11670 -12300
rect 11670 -12370 11740 -12300
rect 11740 -12370 11780 -12300
rect 11780 -12370 11840 -12300
rect 11940 -12370 11960 -12300
rect 11960 -12370 12000 -12300
rect 12000 -12370 12070 -12300
rect 12070 -12370 12110 -12300
rect 12110 -12370 12180 -12300
rect 12270 -12370 12290 -12300
rect 12290 -12370 12330 -12300
rect 12330 -12370 12400 -12300
rect 12400 -12370 12440 -12300
rect 12440 -12370 12510 -12300
rect 11270 -12410 11510 -12370
rect 11600 -12410 11840 -12370
rect 11940 -12410 12180 -12370
rect 12270 -12410 12510 -12370
rect 11270 -12480 11300 -12410
rect 11300 -12480 11340 -12410
rect 11340 -12480 11410 -12410
rect 11410 -12480 11450 -12410
rect 11450 -12480 11510 -12410
rect 11600 -12480 11630 -12410
rect 11630 -12480 11670 -12410
rect 11670 -12480 11740 -12410
rect 11740 -12480 11780 -12410
rect 11780 -12480 11840 -12410
rect 11940 -12480 11960 -12410
rect 11960 -12480 12000 -12410
rect 12000 -12480 12070 -12410
rect 12070 -12480 12110 -12410
rect 12110 -12480 12180 -12410
rect 12270 -12480 12290 -12410
rect 12290 -12480 12330 -12410
rect 12330 -12480 12400 -12410
rect 12400 -12480 12440 -12410
rect 12440 -12480 12510 -12410
rect 19250 -14290 19300 -14230
rect 19300 -14290 19330 -14230
rect 19330 -14290 19400 -14230
rect 19400 -14290 19430 -14230
rect 19430 -14290 19490 -14230
rect 19250 -14320 19490 -14290
rect 19250 -14390 19300 -14320
rect 19300 -14390 19330 -14320
rect 19330 -14390 19400 -14320
rect 19400 -14390 19430 -14320
rect 19430 -14390 19490 -14320
rect 19250 -14420 19490 -14390
rect 19250 -14470 19300 -14420
rect 19300 -14470 19330 -14420
rect 19330 -14470 19400 -14420
rect 19400 -14470 19430 -14420
rect 19430 -14470 19490 -14420
rect 19250 -20360 19300 -20300
rect 19300 -20360 19330 -20300
rect 19330 -20360 19400 -20300
rect 19400 -20360 19430 -20300
rect 19430 -20360 19490 -20300
rect 19250 -20390 19490 -20360
rect 19250 -20460 19300 -20390
rect 19300 -20460 19330 -20390
rect 19330 -20460 19400 -20390
rect 19400 -20460 19430 -20390
rect 19430 -20460 19490 -20390
rect 19250 -20490 19490 -20460
rect 19250 -20540 19300 -20490
rect 19300 -20540 19330 -20490
rect 19330 -20540 19400 -20490
rect 19400 -20540 19430 -20490
rect 19430 -20540 19490 -20490
rect 2390 -22730 2460 -22660
rect 2460 -22730 2500 -22660
rect 2500 -22730 2570 -22660
rect 2570 -22730 2610 -22660
rect 2610 -22730 2630 -22660
rect 2720 -22730 2790 -22660
rect 2790 -22730 2830 -22660
rect 2830 -22730 2900 -22660
rect 2900 -22730 2940 -22660
rect 2940 -22730 2960 -22660
rect 3060 -22730 3120 -22660
rect 3120 -22730 3160 -22660
rect 3160 -22730 3230 -22660
rect 3230 -22730 3270 -22660
rect 3270 -22730 3300 -22660
rect 3390 -22730 3450 -22660
rect 3450 -22730 3490 -22660
rect 3490 -22730 3560 -22660
rect 3560 -22730 3600 -22660
rect 3600 -22730 3630 -22660
rect 2390 -22770 2630 -22730
rect 2720 -22770 2960 -22730
rect 3060 -22770 3300 -22730
rect 3390 -22770 3630 -22730
rect 2390 -22840 2460 -22770
rect 2460 -22840 2500 -22770
rect 2500 -22840 2570 -22770
rect 2570 -22840 2610 -22770
rect 2610 -22840 2630 -22770
rect 2720 -22840 2790 -22770
rect 2790 -22840 2830 -22770
rect 2830 -22840 2900 -22770
rect 2900 -22840 2940 -22770
rect 2940 -22840 2960 -22770
rect 3060 -22840 3120 -22770
rect 3120 -22840 3160 -22770
rect 3160 -22840 3230 -22770
rect 3230 -22840 3270 -22770
rect 3270 -22840 3300 -22770
rect 3390 -22840 3450 -22770
rect 3450 -22840 3490 -22770
rect 3490 -22840 3560 -22770
rect 3560 -22840 3600 -22770
rect 3600 -22840 3630 -22770
rect 2390 -22900 2630 -22840
rect 2720 -22900 2960 -22840
rect 3060 -22900 3300 -22840
rect 3390 -22900 3630 -22840
rect 11270 -22730 11340 -22660
rect 11340 -22730 11380 -22660
rect 11380 -22730 11450 -22660
rect 11450 -22730 11490 -22660
rect 11490 -22730 11510 -22660
rect 11600 -22730 11670 -22660
rect 11670 -22730 11710 -22660
rect 11710 -22730 11780 -22660
rect 11780 -22730 11820 -22660
rect 11820 -22730 11840 -22660
rect 11940 -22730 12000 -22660
rect 12000 -22730 12040 -22660
rect 12040 -22730 12110 -22660
rect 12110 -22730 12150 -22660
rect 12150 -22730 12180 -22660
rect 12270 -22730 12330 -22660
rect 12330 -22730 12370 -22660
rect 12370 -22730 12440 -22660
rect 12440 -22730 12480 -22660
rect 12480 -22730 12510 -22660
rect 11270 -22770 11510 -22730
rect 11600 -22770 11840 -22730
rect 11940 -22770 12180 -22730
rect 12270 -22770 12510 -22730
rect 11270 -22840 11340 -22770
rect 11340 -22840 11380 -22770
rect 11380 -22840 11450 -22770
rect 11450 -22840 11490 -22770
rect 11490 -22840 11510 -22770
rect 11600 -22840 11670 -22770
rect 11670 -22840 11710 -22770
rect 11710 -22840 11780 -22770
rect 11780 -22840 11820 -22770
rect 11820 -22840 11840 -22770
rect 11940 -22840 12000 -22770
rect 12000 -22840 12040 -22770
rect 12040 -22840 12110 -22770
rect 12110 -22840 12150 -22770
rect 12150 -22840 12180 -22770
rect 12270 -22840 12330 -22770
rect 12330 -22840 12370 -22770
rect 12370 -22840 12440 -22770
rect 12440 -22840 12480 -22770
rect 12480 -22840 12510 -22770
rect 11270 -22900 11510 -22840
rect 11600 -22900 11840 -22840
rect 11940 -22900 12180 -22840
rect 12270 -22900 12510 -22840
<< mimcap2 >>
rect -4980 20790 7260 21110
rect -4980 20550 -4670 20790
rect -4430 20550 -4340 20790
rect -4100 20550 -4010 20790
rect -3770 20550 -3680 20790
rect -3440 20550 -3350 20790
rect -3110 20550 -3020 20790
rect -2780 20550 -2690 20790
rect -2450 20550 -2360 20790
rect -2120 20550 -2030 20790
rect -1790 20550 -1700 20790
rect -1460 20550 -1370 20790
rect -1130 20550 -1040 20790
rect -800 20550 -710 20790
rect -470 20550 -380 20790
rect -140 20550 -50 20790
rect 190 20550 280 20790
rect 520 20550 610 20790
rect 850 20550 940 20790
rect 1180 20550 1270 20790
rect 1510 20550 1600 20790
rect 1840 20550 1930 20790
rect 2170 20550 2260 20790
rect 2500 20550 2590 20790
rect 2830 20550 2920 20790
rect 3160 20550 3250 20790
rect 3490 20550 3580 20790
rect 3820 20550 3910 20790
rect 4150 20550 4240 20790
rect 4480 20550 4570 20790
rect 4810 20550 4900 20790
rect 5140 20550 5230 20790
rect 5470 20550 5560 20790
rect 5800 20550 5890 20790
rect 6130 20550 6220 20790
rect 6460 20550 6550 20790
rect 6790 20550 6880 20790
rect 7120 20550 7260 20790
rect -4980 20460 7260 20550
rect -4980 20220 -4670 20460
rect -4430 20220 -4340 20460
rect -4100 20220 -4010 20460
rect -3770 20220 -3680 20460
rect -3440 20220 -3350 20460
rect -3110 20220 -3020 20460
rect -2780 20220 -2690 20460
rect -2450 20220 -2360 20460
rect -2120 20220 -2030 20460
rect -1790 20220 -1700 20460
rect -1460 20220 -1370 20460
rect -1130 20220 -1040 20460
rect -800 20220 -710 20460
rect -470 20220 -380 20460
rect -140 20220 -50 20460
rect 190 20220 280 20460
rect 520 20220 610 20460
rect 850 20220 940 20460
rect 1180 20220 1270 20460
rect 1510 20220 1600 20460
rect 1840 20220 1930 20460
rect 2170 20220 2260 20460
rect 2500 20220 2590 20460
rect 2830 20220 2920 20460
rect 3160 20220 3250 20460
rect 3490 20220 3580 20460
rect 3820 20220 3910 20460
rect 4150 20220 4240 20460
rect 4480 20220 4570 20460
rect 4810 20220 4900 20460
rect 5140 20220 5230 20460
rect 5470 20220 5560 20460
rect 5800 20220 5890 20460
rect 6130 20220 6220 20460
rect 6460 20220 6550 20460
rect 6790 20220 6880 20460
rect 7120 20220 7260 20460
rect -4980 20130 7260 20220
rect -4980 19890 -4670 20130
rect -4430 19890 -4340 20130
rect -4100 19890 -4010 20130
rect -3770 19890 -3680 20130
rect -3440 19890 -3350 20130
rect -3110 19890 -3020 20130
rect -2780 19890 -2690 20130
rect -2450 19890 -2360 20130
rect -2120 19890 -2030 20130
rect -1790 19890 -1700 20130
rect -1460 19890 -1370 20130
rect -1130 19890 -1040 20130
rect -800 19890 -710 20130
rect -470 19890 -380 20130
rect -140 19890 -50 20130
rect 190 19890 280 20130
rect 520 19890 610 20130
rect 850 19890 940 20130
rect 1180 19890 1270 20130
rect 1510 19890 1600 20130
rect 1840 19890 1930 20130
rect 2170 19890 2260 20130
rect 2500 19890 2590 20130
rect 2830 19890 2920 20130
rect 3160 19890 3250 20130
rect 3490 19890 3580 20130
rect 3820 19890 3910 20130
rect 4150 19890 4240 20130
rect 4480 19890 4570 20130
rect 4810 19890 4900 20130
rect 5140 19890 5230 20130
rect 5470 19890 5560 20130
rect 5800 19890 5890 20130
rect 6130 19890 6220 20130
rect 6460 19890 6550 20130
rect 6790 19890 6880 20130
rect 7120 19890 7260 20130
rect -4980 19800 7260 19890
rect -4980 19560 -4670 19800
rect -4430 19560 -4340 19800
rect -4100 19560 -4010 19800
rect -3770 19560 -3680 19800
rect -3440 19560 -3350 19800
rect -3110 19560 -3020 19800
rect -2780 19560 -2690 19800
rect -2450 19560 -2360 19800
rect -2120 19560 -2030 19800
rect -1790 19560 -1700 19800
rect -1460 19560 -1370 19800
rect -1130 19560 -1040 19800
rect -800 19560 -710 19800
rect -470 19560 -380 19800
rect -140 19560 -50 19800
rect 190 19560 280 19800
rect 520 19560 610 19800
rect 850 19560 940 19800
rect 1180 19560 1270 19800
rect 1510 19560 1600 19800
rect 1840 19560 1930 19800
rect 2170 19560 2260 19800
rect 2500 19560 2590 19800
rect 2830 19560 2920 19800
rect 3160 19560 3250 19800
rect 3490 19560 3580 19800
rect 3820 19560 3910 19800
rect 4150 19560 4240 19800
rect 4480 19560 4570 19800
rect 4810 19560 4900 19800
rect 5140 19560 5230 19800
rect 5470 19560 5560 19800
rect 5800 19560 5890 19800
rect 6130 19560 6220 19800
rect 6460 19560 6550 19800
rect 6790 19560 6880 19800
rect 7120 19560 7260 19800
rect -4980 19470 7260 19560
rect -4980 19230 -4670 19470
rect -4430 19230 -4340 19470
rect -4100 19230 -4010 19470
rect -3770 19230 -3680 19470
rect -3440 19230 -3350 19470
rect -3110 19230 -3020 19470
rect -2780 19230 -2690 19470
rect -2450 19230 -2360 19470
rect -2120 19230 -2030 19470
rect -1790 19230 -1700 19470
rect -1460 19230 -1370 19470
rect -1130 19230 -1040 19470
rect -800 19230 -710 19470
rect -470 19230 -380 19470
rect -140 19230 -50 19470
rect 190 19230 280 19470
rect 520 19230 610 19470
rect 850 19230 940 19470
rect 1180 19230 1270 19470
rect 1510 19230 1600 19470
rect 1840 19230 1930 19470
rect 2170 19230 2260 19470
rect 2500 19230 2590 19470
rect 2830 19230 2920 19470
rect 3160 19230 3250 19470
rect 3490 19230 3580 19470
rect 3820 19230 3910 19470
rect 4150 19230 4240 19470
rect 4480 19230 4570 19470
rect 4810 19230 4900 19470
rect 5140 19230 5230 19470
rect 5470 19230 5560 19470
rect 5800 19230 5890 19470
rect 6130 19230 6220 19470
rect 6460 19230 6550 19470
rect 6790 19230 6880 19470
rect 7120 19230 7260 19470
rect -4980 19140 7260 19230
rect -4980 18900 -4670 19140
rect -4430 18900 -4340 19140
rect -4100 18900 -4010 19140
rect -3770 18900 -3680 19140
rect -3440 18900 -3350 19140
rect -3110 18900 -3020 19140
rect -2780 18900 -2690 19140
rect -2450 18900 -2360 19140
rect -2120 18900 -2030 19140
rect -1790 18900 -1700 19140
rect -1460 18900 -1370 19140
rect -1130 18900 -1040 19140
rect -800 18900 -710 19140
rect -470 18900 -380 19140
rect -140 18900 -50 19140
rect 190 18900 280 19140
rect 520 18900 610 19140
rect 850 18900 940 19140
rect 1180 18900 1270 19140
rect 1510 18900 1600 19140
rect 1840 18900 1930 19140
rect 2170 18900 2260 19140
rect 2500 18900 2590 19140
rect 2830 18900 2920 19140
rect 3160 18900 3250 19140
rect 3490 18900 3580 19140
rect 3820 18900 3910 19140
rect 4150 18900 4240 19140
rect 4480 18900 4570 19140
rect 4810 18900 4900 19140
rect 5140 18900 5230 19140
rect 5470 18900 5560 19140
rect 5800 18900 5890 19140
rect 6130 18900 6220 19140
rect 6460 18900 6550 19140
rect 6790 18900 6880 19140
rect 7120 18900 7260 19140
rect -4980 18810 7260 18900
rect -4980 18570 -4670 18810
rect -4430 18570 -4340 18810
rect -4100 18570 -4010 18810
rect -3770 18570 -3680 18810
rect -3440 18570 -3350 18810
rect -3110 18570 -3020 18810
rect -2780 18570 -2690 18810
rect -2450 18570 -2360 18810
rect -2120 18570 -2030 18810
rect -1790 18570 -1700 18810
rect -1460 18570 -1370 18810
rect -1130 18570 -1040 18810
rect -800 18570 -710 18810
rect -470 18570 -380 18810
rect -140 18570 -50 18810
rect 190 18570 280 18810
rect 520 18570 610 18810
rect 850 18570 940 18810
rect 1180 18570 1270 18810
rect 1510 18570 1600 18810
rect 1840 18570 1930 18810
rect 2170 18570 2260 18810
rect 2500 18570 2590 18810
rect 2830 18570 2920 18810
rect 3160 18570 3250 18810
rect 3490 18570 3580 18810
rect 3820 18570 3910 18810
rect 4150 18570 4240 18810
rect 4480 18570 4570 18810
rect 4810 18570 4900 18810
rect 5140 18570 5230 18810
rect 5470 18570 5560 18810
rect 5800 18570 5890 18810
rect 6130 18570 6220 18810
rect 6460 18570 6550 18810
rect 6790 18570 6880 18810
rect 7120 18570 7260 18810
rect -4980 18480 7260 18570
rect -4980 18240 -4670 18480
rect -4430 18240 -4340 18480
rect -4100 18240 -4010 18480
rect -3770 18240 -3680 18480
rect -3440 18240 -3350 18480
rect -3110 18240 -3020 18480
rect -2780 18240 -2690 18480
rect -2450 18240 -2360 18480
rect -2120 18240 -2030 18480
rect -1790 18240 -1700 18480
rect -1460 18240 -1370 18480
rect -1130 18240 -1040 18480
rect -800 18240 -710 18480
rect -470 18240 -380 18480
rect -140 18240 -50 18480
rect 190 18240 280 18480
rect 520 18240 610 18480
rect 850 18240 940 18480
rect 1180 18240 1270 18480
rect 1510 18240 1600 18480
rect 1840 18240 1930 18480
rect 2170 18240 2260 18480
rect 2500 18240 2590 18480
rect 2830 18240 2920 18480
rect 3160 18240 3250 18480
rect 3490 18240 3580 18480
rect 3820 18240 3910 18480
rect 4150 18240 4240 18480
rect 4480 18240 4570 18480
rect 4810 18240 4900 18480
rect 5140 18240 5230 18480
rect 5470 18240 5560 18480
rect 5800 18240 5890 18480
rect 6130 18240 6220 18480
rect 6460 18240 6550 18480
rect 6790 18240 6880 18480
rect 7120 18240 7260 18480
rect -4980 18150 7260 18240
rect -4980 17910 -4670 18150
rect -4430 17910 -4340 18150
rect -4100 17910 -4010 18150
rect -3770 17910 -3680 18150
rect -3440 17910 -3350 18150
rect -3110 17910 -3020 18150
rect -2780 17910 -2690 18150
rect -2450 17910 -2360 18150
rect -2120 17910 -2030 18150
rect -1790 17910 -1700 18150
rect -1460 17910 -1370 18150
rect -1130 17910 -1040 18150
rect -800 17910 -710 18150
rect -470 17910 -380 18150
rect -140 17910 -50 18150
rect 190 17910 280 18150
rect 520 17910 610 18150
rect 850 17910 940 18150
rect 1180 17910 1270 18150
rect 1510 17910 1600 18150
rect 1840 17910 1930 18150
rect 2170 17910 2260 18150
rect 2500 17910 2590 18150
rect 2830 17910 2920 18150
rect 3160 17910 3250 18150
rect 3490 17910 3580 18150
rect 3820 17910 3910 18150
rect 4150 17910 4240 18150
rect 4480 17910 4570 18150
rect 4810 17910 4900 18150
rect 5140 17910 5230 18150
rect 5470 17910 5560 18150
rect 5800 17910 5890 18150
rect 6130 17910 6220 18150
rect 6460 17910 6550 18150
rect 6790 17910 6880 18150
rect 7120 17910 7260 18150
rect -4980 17820 7260 17910
rect -4980 17580 -4670 17820
rect -4430 17580 -4340 17820
rect -4100 17580 -4010 17820
rect -3770 17580 -3680 17820
rect -3440 17580 -3350 17820
rect -3110 17580 -3020 17820
rect -2780 17580 -2690 17820
rect -2450 17580 -2360 17820
rect -2120 17580 -2030 17820
rect -1790 17580 -1700 17820
rect -1460 17580 -1370 17820
rect -1130 17580 -1040 17820
rect -800 17580 -710 17820
rect -470 17580 -380 17820
rect -140 17580 -50 17820
rect 190 17580 280 17820
rect 520 17580 610 17820
rect 850 17580 940 17820
rect 1180 17580 1270 17820
rect 1510 17580 1600 17820
rect 1840 17580 1930 17820
rect 2170 17580 2260 17820
rect 2500 17580 2590 17820
rect 2830 17580 2920 17820
rect 3160 17580 3250 17820
rect 3490 17580 3580 17820
rect 3820 17580 3910 17820
rect 4150 17580 4240 17820
rect 4480 17580 4570 17820
rect 4810 17580 4900 17820
rect 5140 17580 5230 17820
rect 5470 17580 5560 17820
rect 5800 17580 5890 17820
rect 6130 17580 6220 17820
rect 6460 17580 6550 17820
rect 6790 17580 6880 17820
rect 7120 17580 7260 17820
rect -4980 17490 7260 17580
rect -4980 17250 -4670 17490
rect -4430 17250 -4340 17490
rect -4100 17250 -4010 17490
rect -3770 17250 -3680 17490
rect -3440 17250 -3350 17490
rect -3110 17250 -3020 17490
rect -2780 17250 -2690 17490
rect -2450 17250 -2360 17490
rect -2120 17250 -2030 17490
rect -1790 17250 -1700 17490
rect -1460 17250 -1370 17490
rect -1130 17250 -1040 17490
rect -800 17250 -710 17490
rect -470 17250 -380 17490
rect -140 17250 -50 17490
rect 190 17250 280 17490
rect 520 17250 610 17490
rect 850 17250 940 17490
rect 1180 17250 1270 17490
rect 1510 17250 1600 17490
rect 1840 17250 1930 17490
rect 2170 17250 2260 17490
rect 2500 17250 2590 17490
rect 2830 17250 2920 17490
rect 3160 17250 3250 17490
rect 3490 17250 3580 17490
rect 3820 17250 3910 17490
rect 4150 17250 4240 17490
rect 4480 17250 4570 17490
rect 4810 17250 4900 17490
rect 5140 17250 5230 17490
rect 5470 17250 5560 17490
rect 5800 17250 5890 17490
rect 6130 17250 6220 17490
rect 6460 17250 6550 17490
rect 6790 17250 6880 17490
rect 7120 17250 7260 17490
rect -4980 17160 7260 17250
rect -4980 16920 -4670 17160
rect -4430 16920 -4340 17160
rect -4100 16920 -4010 17160
rect -3770 16920 -3680 17160
rect -3440 16920 -3350 17160
rect -3110 16920 -3020 17160
rect -2780 16920 -2690 17160
rect -2450 16920 -2360 17160
rect -2120 16920 -2030 17160
rect -1790 16920 -1700 17160
rect -1460 16920 -1370 17160
rect -1130 16920 -1040 17160
rect -800 16920 -710 17160
rect -470 16920 -380 17160
rect -140 16920 -50 17160
rect 190 16920 280 17160
rect 520 16920 610 17160
rect 850 16920 940 17160
rect 1180 16920 1270 17160
rect 1510 16920 1600 17160
rect 1840 16920 1930 17160
rect 2170 16920 2260 17160
rect 2500 16920 2590 17160
rect 2830 16920 2920 17160
rect 3160 16920 3250 17160
rect 3490 16920 3580 17160
rect 3820 16920 3910 17160
rect 4150 16920 4240 17160
rect 4480 16920 4570 17160
rect 4810 16920 4900 17160
rect 5140 16920 5230 17160
rect 5470 16920 5560 17160
rect 5800 16920 5890 17160
rect 6130 16920 6220 17160
rect 6460 16920 6550 17160
rect 6790 16920 6880 17160
rect 7120 16920 7260 17160
rect -4980 16830 7260 16920
rect -4980 16590 -4670 16830
rect -4430 16590 -4340 16830
rect -4100 16590 -4010 16830
rect -3770 16590 -3680 16830
rect -3440 16590 -3350 16830
rect -3110 16590 -3020 16830
rect -2780 16590 -2690 16830
rect -2450 16590 -2360 16830
rect -2120 16590 -2030 16830
rect -1790 16590 -1700 16830
rect -1460 16590 -1370 16830
rect -1130 16590 -1040 16830
rect -800 16590 -710 16830
rect -470 16590 -380 16830
rect -140 16590 -50 16830
rect 190 16590 280 16830
rect 520 16590 610 16830
rect 850 16590 940 16830
rect 1180 16590 1270 16830
rect 1510 16590 1600 16830
rect 1840 16590 1930 16830
rect 2170 16590 2260 16830
rect 2500 16590 2590 16830
rect 2830 16590 2920 16830
rect 3160 16590 3250 16830
rect 3490 16590 3580 16830
rect 3820 16590 3910 16830
rect 4150 16590 4240 16830
rect 4480 16590 4570 16830
rect 4810 16590 4900 16830
rect 5140 16590 5230 16830
rect 5470 16590 5560 16830
rect 5800 16590 5890 16830
rect 6130 16590 6220 16830
rect 6460 16590 6550 16830
rect 6790 16590 6880 16830
rect 7120 16590 7260 16830
rect -4980 16500 7260 16590
rect -4980 16260 -4670 16500
rect -4430 16260 -4340 16500
rect -4100 16260 -4010 16500
rect -3770 16260 -3680 16500
rect -3440 16260 -3350 16500
rect -3110 16260 -3020 16500
rect -2780 16260 -2690 16500
rect -2450 16260 -2360 16500
rect -2120 16260 -2030 16500
rect -1790 16260 -1700 16500
rect -1460 16260 -1370 16500
rect -1130 16260 -1040 16500
rect -800 16260 -710 16500
rect -470 16260 -380 16500
rect -140 16260 -50 16500
rect 190 16260 280 16500
rect 520 16260 610 16500
rect 850 16260 940 16500
rect 1180 16260 1270 16500
rect 1510 16260 1600 16500
rect 1840 16260 1930 16500
rect 2170 16260 2260 16500
rect 2500 16260 2590 16500
rect 2830 16260 2920 16500
rect 3160 16260 3250 16500
rect 3490 16260 3580 16500
rect 3820 16260 3910 16500
rect 4150 16260 4240 16500
rect 4480 16260 4570 16500
rect 4810 16260 4900 16500
rect 5140 16260 5230 16500
rect 5470 16260 5560 16500
rect 5800 16260 5890 16500
rect 6130 16260 6220 16500
rect 6460 16260 6550 16500
rect 6790 16260 6880 16500
rect 7120 16260 7260 16500
rect -4980 16170 7260 16260
rect -4980 15930 -4670 16170
rect -4430 15930 -4340 16170
rect -4100 15930 -4010 16170
rect -3770 15930 -3680 16170
rect -3440 15930 -3350 16170
rect -3110 15930 -3020 16170
rect -2780 15930 -2690 16170
rect -2450 15930 -2360 16170
rect -2120 15930 -2030 16170
rect -1790 15930 -1700 16170
rect -1460 15930 -1370 16170
rect -1130 15930 -1040 16170
rect -800 15930 -710 16170
rect -470 15930 -380 16170
rect -140 15930 -50 16170
rect 190 15930 280 16170
rect 520 15930 610 16170
rect 850 15930 940 16170
rect 1180 15930 1270 16170
rect 1510 15930 1600 16170
rect 1840 15930 1930 16170
rect 2170 15930 2260 16170
rect 2500 15930 2590 16170
rect 2830 15930 2920 16170
rect 3160 15930 3250 16170
rect 3490 15930 3580 16170
rect 3820 15930 3910 16170
rect 4150 15930 4240 16170
rect 4480 15930 4570 16170
rect 4810 15930 4900 16170
rect 5140 15930 5230 16170
rect 5470 15930 5560 16170
rect 5800 15930 5890 16170
rect 6130 15930 6220 16170
rect 6460 15930 6550 16170
rect 6790 15930 6880 16170
rect 7120 15930 7260 16170
rect -4980 15840 7260 15930
rect -4980 15600 -4670 15840
rect -4430 15600 -4340 15840
rect -4100 15600 -4010 15840
rect -3770 15600 -3680 15840
rect -3440 15600 -3350 15840
rect -3110 15600 -3020 15840
rect -2780 15600 -2690 15840
rect -2450 15600 -2360 15840
rect -2120 15600 -2030 15840
rect -1790 15600 -1700 15840
rect -1460 15600 -1370 15840
rect -1130 15600 -1040 15840
rect -800 15600 -710 15840
rect -470 15600 -380 15840
rect -140 15600 -50 15840
rect 190 15600 280 15840
rect 520 15600 610 15840
rect 850 15600 940 15840
rect 1180 15600 1270 15840
rect 1510 15600 1600 15840
rect 1840 15600 1930 15840
rect 2170 15600 2260 15840
rect 2500 15600 2590 15840
rect 2830 15600 2920 15840
rect 3160 15600 3250 15840
rect 3490 15600 3580 15840
rect 3820 15600 3910 15840
rect 4150 15600 4240 15840
rect 4480 15600 4570 15840
rect 4810 15600 4900 15840
rect 5140 15600 5230 15840
rect 5470 15600 5560 15840
rect 5800 15600 5890 15840
rect 6130 15600 6220 15840
rect 6460 15600 6550 15840
rect 6790 15600 6880 15840
rect 7120 15600 7260 15840
rect -4980 15510 7260 15600
rect -4980 15270 -4670 15510
rect -4430 15270 -4340 15510
rect -4100 15270 -4010 15510
rect -3770 15270 -3680 15510
rect -3440 15270 -3350 15510
rect -3110 15270 -3020 15510
rect -2780 15270 -2690 15510
rect -2450 15270 -2360 15510
rect -2120 15270 -2030 15510
rect -1790 15270 -1700 15510
rect -1460 15270 -1370 15510
rect -1130 15270 -1040 15510
rect -800 15270 -710 15510
rect -470 15270 -380 15510
rect -140 15270 -50 15510
rect 190 15270 280 15510
rect 520 15270 610 15510
rect 850 15270 940 15510
rect 1180 15270 1270 15510
rect 1510 15270 1600 15510
rect 1840 15270 1930 15510
rect 2170 15270 2260 15510
rect 2500 15270 2590 15510
rect 2830 15270 2920 15510
rect 3160 15270 3250 15510
rect 3490 15270 3580 15510
rect 3820 15270 3910 15510
rect 4150 15270 4240 15510
rect 4480 15270 4570 15510
rect 4810 15270 4900 15510
rect 5140 15270 5230 15510
rect 5470 15270 5560 15510
rect 5800 15270 5890 15510
rect 6130 15270 6220 15510
rect 6460 15270 6550 15510
rect 6790 15270 6880 15510
rect 7120 15270 7260 15510
rect -4980 15180 7260 15270
rect -4980 14940 -4670 15180
rect -4430 14940 -4340 15180
rect -4100 14940 -4010 15180
rect -3770 14940 -3680 15180
rect -3440 14940 -3350 15180
rect -3110 14940 -3020 15180
rect -2780 14940 -2690 15180
rect -2450 14940 -2360 15180
rect -2120 14940 -2030 15180
rect -1790 14940 -1700 15180
rect -1460 14940 -1370 15180
rect -1130 14940 -1040 15180
rect -800 14940 -710 15180
rect -470 14940 -380 15180
rect -140 14940 -50 15180
rect 190 14940 280 15180
rect 520 14940 610 15180
rect 850 14940 940 15180
rect 1180 14940 1270 15180
rect 1510 14940 1600 15180
rect 1840 14940 1930 15180
rect 2170 14940 2260 15180
rect 2500 14940 2590 15180
rect 2830 14940 2920 15180
rect 3160 14940 3250 15180
rect 3490 14940 3580 15180
rect 3820 14940 3910 15180
rect 4150 14940 4240 15180
rect 4480 14940 4570 15180
rect 4810 14940 4900 15180
rect 5140 14940 5230 15180
rect 5470 14940 5560 15180
rect 5800 14940 5890 15180
rect 6130 14940 6220 15180
rect 6460 14940 6550 15180
rect 6790 14940 6880 15180
rect 7120 14940 7260 15180
rect -4980 14850 7260 14940
rect -4980 14610 -4670 14850
rect -4430 14610 -4340 14850
rect -4100 14610 -4010 14850
rect -3770 14610 -3680 14850
rect -3440 14610 -3350 14850
rect -3110 14610 -3020 14850
rect -2780 14610 -2690 14850
rect -2450 14610 -2360 14850
rect -2120 14610 -2030 14850
rect -1790 14610 -1700 14850
rect -1460 14610 -1370 14850
rect -1130 14610 -1040 14850
rect -800 14610 -710 14850
rect -470 14610 -380 14850
rect -140 14610 -50 14850
rect 190 14610 280 14850
rect 520 14610 610 14850
rect 850 14610 940 14850
rect 1180 14610 1270 14850
rect 1510 14610 1600 14850
rect 1840 14610 1930 14850
rect 2170 14610 2260 14850
rect 2500 14610 2590 14850
rect 2830 14610 2920 14850
rect 3160 14610 3250 14850
rect 3490 14610 3580 14850
rect 3820 14610 3910 14850
rect 4150 14610 4240 14850
rect 4480 14610 4570 14850
rect 4810 14610 4900 14850
rect 5140 14610 5230 14850
rect 5470 14610 5560 14850
rect 5800 14610 5890 14850
rect 6130 14610 6220 14850
rect 6460 14610 6550 14850
rect 6790 14610 6880 14850
rect 7120 14610 7260 14850
rect -4980 14520 7260 14610
rect -4980 14280 -4670 14520
rect -4430 14280 -4340 14520
rect -4100 14280 -4010 14520
rect -3770 14280 -3680 14520
rect -3440 14280 -3350 14520
rect -3110 14280 -3020 14520
rect -2780 14280 -2690 14520
rect -2450 14280 -2360 14520
rect -2120 14280 -2030 14520
rect -1790 14280 -1700 14520
rect -1460 14280 -1370 14520
rect -1130 14280 -1040 14520
rect -800 14280 -710 14520
rect -470 14280 -380 14520
rect -140 14280 -50 14520
rect 190 14280 280 14520
rect 520 14280 610 14520
rect 850 14280 940 14520
rect 1180 14280 1270 14520
rect 1510 14280 1600 14520
rect 1840 14280 1930 14520
rect 2170 14280 2260 14520
rect 2500 14280 2590 14520
rect 2830 14280 2920 14520
rect 3160 14280 3250 14520
rect 3490 14280 3580 14520
rect 3820 14280 3910 14520
rect 4150 14280 4240 14520
rect 4480 14280 4570 14520
rect 4810 14280 4900 14520
rect 5140 14280 5230 14520
rect 5470 14280 5560 14520
rect 5800 14280 5890 14520
rect 6130 14280 6220 14520
rect 6460 14280 6550 14520
rect 6790 14280 6880 14520
rect 7120 14280 7260 14520
rect -4980 14190 7260 14280
rect -4980 13950 -4670 14190
rect -4430 13950 -4340 14190
rect -4100 13950 -4010 14190
rect -3770 13950 -3680 14190
rect -3440 13950 -3350 14190
rect -3110 13950 -3020 14190
rect -2780 13950 -2690 14190
rect -2450 13950 -2360 14190
rect -2120 13950 -2030 14190
rect -1790 13950 -1700 14190
rect -1460 13950 -1370 14190
rect -1130 13950 -1040 14190
rect -800 13950 -710 14190
rect -470 13950 -380 14190
rect -140 13950 -50 14190
rect 190 13950 280 14190
rect 520 13950 610 14190
rect 850 13950 940 14190
rect 1180 13950 1270 14190
rect 1510 13950 1600 14190
rect 1840 13950 1930 14190
rect 2170 13950 2260 14190
rect 2500 13950 2590 14190
rect 2830 13950 2920 14190
rect 3160 13950 3250 14190
rect 3490 13950 3580 14190
rect 3820 13950 3910 14190
rect 4150 13950 4240 14190
rect 4480 13950 4570 14190
rect 4810 13950 4900 14190
rect 5140 13950 5230 14190
rect 5470 13950 5560 14190
rect 5800 13950 5890 14190
rect 6130 13950 6220 14190
rect 6460 13950 6550 14190
rect 6790 13950 6880 14190
rect 7120 13950 7260 14190
rect -4980 13860 7260 13950
rect -4980 13620 -4670 13860
rect -4430 13620 -4340 13860
rect -4100 13620 -4010 13860
rect -3770 13620 -3680 13860
rect -3440 13620 -3350 13860
rect -3110 13620 -3020 13860
rect -2780 13620 -2690 13860
rect -2450 13620 -2360 13860
rect -2120 13620 -2030 13860
rect -1790 13620 -1700 13860
rect -1460 13620 -1370 13860
rect -1130 13620 -1040 13860
rect -800 13620 -710 13860
rect -470 13620 -380 13860
rect -140 13620 -50 13860
rect 190 13620 280 13860
rect 520 13620 610 13860
rect 850 13620 940 13860
rect 1180 13620 1270 13860
rect 1510 13620 1600 13860
rect 1840 13620 1930 13860
rect 2170 13620 2260 13860
rect 2500 13620 2590 13860
rect 2830 13620 2920 13860
rect 3160 13620 3250 13860
rect 3490 13620 3580 13860
rect 3820 13620 3910 13860
rect 4150 13620 4240 13860
rect 4480 13620 4570 13860
rect 4810 13620 4900 13860
rect 5140 13620 5230 13860
rect 5470 13620 5560 13860
rect 5800 13620 5890 13860
rect 6130 13620 6220 13860
rect 6460 13620 6550 13860
rect 6790 13620 6880 13860
rect 7120 13620 7260 13860
rect -4980 13530 7260 13620
rect -4980 13290 -4670 13530
rect -4430 13290 -4340 13530
rect -4100 13290 -4010 13530
rect -3770 13290 -3680 13530
rect -3440 13290 -3350 13530
rect -3110 13290 -3020 13530
rect -2780 13290 -2690 13530
rect -2450 13290 -2360 13530
rect -2120 13290 -2030 13530
rect -1790 13290 -1700 13530
rect -1460 13290 -1370 13530
rect -1130 13290 -1040 13530
rect -800 13290 -710 13530
rect -470 13290 -380 13530
rect -140 13290 -50 13530
rect 190 13290 280 13530
rect 520 13290 610 13530
rect 850 13290 940 13530
rect 1180 13290 1270 13530
rect 1510 13290 1600 13530
rect 1840 13290 1930 13530
rect 2170 13290 2260 13530
rect 2500 13290 2590 13530
rect 2830 13290 2920 13530
rect 3160 13290 3250 13530
rect 3490 13290 3580 13530
rect 3820 13290 3910 13530
rect 4150 13290 4240 13530
rect 4480 13290 4570 13530
rect 4810 13290 4900 13530
rect 5140 13290 5230 13530
rect 5470 13290 5560 13530
rect 5800 13290 5890 13530
rect 6130 13290 6220 13530
rect 6460 13290 6550 13530
rect 6790 13290 6880 13530
rect 7120 13290 7260 13530
rect -4980 13200 7260 13290
rect -4980 12960 -4670 13200
rect -4430 12960 -4340 13200
rect -4100 12960 -4010 13200
rect -3770 12960 -3680 13200
rect -3440 12960 -3350 13200
rect -3110 12960 -3020 13200
rect -2780 12960 -2690 13200
rect -2450 12960 -2360 13200
rect -2120 12960 -2030 13200
rect -1790 12960 -1700 13200
rect -1460 12960 -1370 13200
rect -1130 12960 -1040 13200
rect -800 12960 -710 13200
rect -470 12960 -380 13200
rect -140 12960 -50 13200
rect 190 12960 280 13200
rect 520 12960 610 13200
rect 850 12960 940 13200
rect 1180 12960 1270 13200
rect 1510 12960 1600 13200
rect 1840 12960 1930 13200
rect 2170 12960 2260 13200
rect 2500 12960 2590 13200
rect 2830 12960 2920 13200
rect 3160 12960 3250 13200
rect 3490 12960 3580 13200
rect 3820 12960 3910 13200
rect 4150 12960 4240 13200
rect 4480 12960 4570 13200
rect 4810 12960 4900 13200
rect 5140 12960 5230 13200
rect 5470 12960 5560 13200
rect 5800 12960 5890 13200
rect 6130 12960 6220 13200
rect 6460 12960 6550 13200
rect 6790 12960 6880 13200
rect 7120 12960 7260 13200
rect -4980 12870 7260 12960
rect -4980 12630 -4670 12870
rect -4430 12630 -4340 12870
rect -4100 12630 -4010 12870
rect -3770 12630 -3680 12870
rect -3440 12630 -3350 12870
rect -3110 12630 -3020 12870
rect -2780 12630 -2690 12870
rect -2450 12630 -2360 12870
rect -2120 12630 -2030 12870
rect -1790 12630 -1700 12870
rect -1460 12630 -1370 12870
rect -1130 12630 -1040 12870
rect -800 12630 -710 12870
rect -470 12630 -380 12870
rect -140 12630 -50 12870
rect 190 12630 280 12870
rect 520 12630 610 12870
rect 850 12630 940 12870
rect 1180 12630 1270 12870
rect 1510 12630 1600 12870
rect 1840 12630 1930 12870
rect 2170 12630 2260 12870
rect 2500 12630 2590 12870
rect 2830 12630 2920 12870
rect 3160 12630 3250 12870
rect 3490 12630 3580 12870
rect 3820 12630 3910 12870
rect 4150 12630 4240 12870
rect 4480 12630 4570 12870
rect 4810 12630 4900 12870
rect 5140 12630 5230 12870
rect 5470 12630 5560 12870
rect 5800 12630 5890 12870
rect 6130 12630 6220 12870
rect 6460 12630 6550 12870
rect 6790 12630 6880 12870
rect 7120 12630 7260 12870
rect -4980 12540 7260 12630
rect -4980 12300 -4670 12540
rect -4430 12300 -4340 12540
rect -4100 12300 -4010 12540
rect -3770 12300 -3680 12540
rect -3440 12300 -3350 12540
rect -3110 12300 -3020 12540
rect -2780 12300 -2690 12540
rect -2450 12300 -2360 12540
rect -2120 12300 -2030 12540
rect -1790 12300 -1700 12540
rect -1460 12300 -1370 12540
rect -1130 12300 -1040 12540
rect -800 12300 -710 12540
rect -470 12300 -380 12540
rect -140 12300 -50 12540
rect 190 12300 280 12540
rect 520 12300 610 12540
rect 850 12300 940 12540
rect 1180 12300 1270 12540
rect 1510 12300 1600 12540
rect 1840 12300 1930 12540
rect 2170 12300 2260 12540
rect 2500 12300 2590 12540
rect 2830 12300 2920 12540
rect 3160 12300 3250 12540
rect 3490 12300 3580 12540
rect 3820 12300 3910 12540
rect 4150 12300 4240 12540
rect 4480 12300 4570 12540
rect 4810 12300 4900 12540
rect 5140 12300 5230 12540
rect 5470 12300 5560 12540
rect 5800 12300 5890 12540
rect 6130 12300 6220 12540
rect 6460 12300 6550 12540
rect 6790 12300 6880 12540
rect 7120 12300 7260 12540
rect -4980 12210 7260 12300
rect -4980 11970 -4670 12210
rect -4430 11970 -4340 12210
rect -4100 11970 -4010 12210
rect -3770 11970 -3680 12210
rect -3440 11970 -3350 12210
rect -3110 11970 -3020 12210
rect -2780 11970 -2690 12210
rect -2450 11970 -2360 12210
rect -2120 11970 -2030 12210
rect -1790 11970 -1700 12210
rect -1460 11970 -1370 12210
rect -1130 11970 -1040 12210
rect -800 11970 -710 12210
rect -470 11970 -380 12210
rect -140 11970 -50 12210
rect 190 11970 280 12210
rect 520 11970 610 12210
rect 850 11970 940 12210
rect 1180 11970 1270 12210
rect 1510 11970 1600 12210
rect 1840 11970 1930 12210
rect 2170 11970 2260 12210
rect 2500 11970 2590 12210
rect 2830 11970 2920 12210
rect 3160 11970 3250 12210
rect 3490 11970 3580 12210
rect 3820 11970 3910 12210
rect 4150 11970 4240 12210
rect 4480 11970 4570 12210
rect 4810 11970 4900 12210
rect 5140 11970 5230 12210
rect 5470 11970 5560 12210
rect 5800 11970 5890 12210
rect 6130 11970 6220 12210
rect 6460 11970 6550 12210
rect 6790 11970 6880 12210
rect 7120 11970 7260 12210
rect -4980 11880 7260 11970
rect -4980 11640 -4670 11880
rect -4430 11640 -4340 11880
rect -4100 11640 -4010 11880
rect -3770 11640 -3680 11880
rect -3440 11640 -3350 11880
rect -3110 11640 -3020 11880
rect -2780 11640 -2690 11880
rect -2450 11640 -2360 11880
rect -2120 11640 -2030 11880
rect -1790 11640 -1700 11880
rect -1460 11640 -1370 11880
rect -1130 11640 -1040 11880
rect -800 11640 -710 11880
rect -470 11640 -380 11880
rect -140 11640 -50 11880
rect 190 11640 280 11880
rect 520 11640 610 11880
rect 850 11640 940 11880
rect 1180 11640 1270 11880
rect 1510 11640 1600 11880
rect 1840 11640 1930 11880
rect 2170 11640 2260 11880
rect 2500 11640 2590 11880
rect 2830 11640 2920 11880
rect 3160 11640 3250 11880
rect 3490 11640 3580 11880
rect 3820 11640 3910 11880
rect 4150 11640 4240 11880
rect 4480 11640 4570 11880
rect 4810 11640 4900 11880
rect 5140 11640 5230 11880
rect 5470 11640 5560 11880
rect 5800 11640 5890 11880
rect 6130 11640 6220 11880
rect 6460 11640 6550 11880
rect 6790 11640 6880 11880
rect 7120 11640 7260 11880
rect -4980 11550 7260 11640
rect -4980 11310 -4670 11550
rect -4430 11310 -4340 11550
rect -4100 11310 -4010 11550
rect -3770 11310 -3680 11550
rect -3440 11310 -3350 11550
rect -3110 11310 -3020 11550
rect -2780 11310 -2690 11550
rect -2450 11310 -2360 11550
rect -2120 11310 -2030 11550
rect -1790 11310 -1700 11550
rect -1460 11310 -1370 11550
rect -1130 11310 -1040 11550
rect -800 11310 -710 11550
rect -470 11310 -380 11550
rect -140 11310 -50 11550
rect 190 11310 280 11550
rect 520 11310 610 11550
rect 850 11310 940 11550
rect 1180 11310 1270 11550
rect 1510 11310 1600 11550
rect 1840 11310 1930 11550
rect 2170 11310 2260 11550
rect 2500 11310 2590 11550
rect 2830 11310 2920 11550
rect 3160 11310 3250 11550
rect 3490 11310 3580 11550
rect 3820 11310 3910 11550
rect 4150 11310 4240 11550
rect 4480 11310 4570 11550
rect 4810 11310 4900 11550
rect 5140 11310 5230 11550
rect 5470 11310 5560 11550
rect 5800 11310 5890 11550
rect 6130 11310 6220 11550
rect 6460 11310 6550 11550
rect 6790 11310 6880 11550
rect 7120 11310 7260 11550
rect -4980 11220 7260 11310
rect -4980 10980 -4670 11220
rect -4430 10980 -4340 11220
rect -4100 10980 -4010 11220
rect -3770 10980 -3680 11220
rect -3440 10980 -3350 11220
rect -3110 10980 -3020 11220
rect -2780 10980 -2690 11220
rect -2450 10980 -2360 11220
rect -2120 10980 -2030 11220
rect -1790 10980 -1700 11220
rect -1460 10980 -1370 11220
rect -1130 10980 -1040 11220
rect -800 10980 -710 11220
rect -470 10980 -380 11220
rect -140 10980 -50 11220
rect 190 10980 280 11220
rect 520 10980 610 11220
rect 850 10980 940 11220
rect 1180 10980 1270 11220
rect 1510 10980 1600 11220
rect 1840 10980 1930 11220
rect 2170 10980 2260 11220
rect 2500 10980 2590 11220
rect 2830 10980 2920 11220
rect 3160 10980 3250 11220
rect 3490 10980 3580 11220
rect 3820 10980 3910 11220
rect 4150 10980 4240 11220
rect 4480 10980 4570 11220
rect 4810 10980 4900 11220
rect 5140 10980 5230 11220
rect 5470 10980 5560 11220
rect 5800 10980 5890 11220
rect 6130 10980 6220 11220
rect 6460 10980 6550 11220
rect 6790 10980 6880 11220
rect 7120 10980 7260 11220
rect -4980 10890 7260 10980
rect -4980 10650 -4670 10890
rect -4430 10650 -4340 10890
rect -4100 10650 -4010 10890
rect -3770 10650 -3680 10890
rect -3440 10650 -3350 10890
rect -3110 10650 -3020 10890
rect -2780 10650 -2690 10890
rect -2450 10650 -2360 10890
rect -2120 10650 -2030 10890
rect -1790 10650 -1700 10890
rect -1460 10650 -1370 10890
rect -1130 10650 -1040 10890
rect -800 10650 -710 10890
rect -470 10650 -380 10890
rect -140 10650 -50 10890
rect 190 10650 280 10890
rect 520 10650 610 10890
rect 850 10650 940 10890
rect 1180 10650 1270 10890
rect 1510 10650 1600 10890
rect 1840 10650 1930 10890
rect 2170 10650 2260 10890
rect 2500 10650 2590 10890
rect 2830 10650 2920 10890
rect 3160 10650 3250 10890
rect 3490 10650 3580 10890
rect 3820 10650 3910 10890
rect 4150 10650 4240 10890
rect 4480 10650 4570 10890
rect 4810 10650 4900 10890
rect 5140 10650 5230 10890
rect 5470 10650 5560 10890
rect 5800 10650 5890 10890
rect 6130 10650 6220 10890
rect 6460 10650 6550 10890
rect 6790 10650 6880 10890
rect 7120 10650 7260 10890
rect -4980 10560 7260 10650
rect -4980 10320 -4670 10560
rect -4430 10320 -4340 10560
rect -4100 10320 -4010 10560
rect -3770 10320 -3680 10560
rect -3440 10320 -3350 10560
rect -3110 10320 -3020 10560
rect -2780 10320 -2690 10560
rect -2450 10320 -2360 10560
rect -2120 10320 -2030 10560
rect -1790 10320 -1700 10560
rect -1460 10320 -1370 10560
rect -1130 10320 -1040 10560
rect -800 10320 -710 10560
rect -470 10320 -380 10560
rect -140 10320 -50 10560
rect 190 10320 280 10560
rect 520 10320 610 10560
rect 850 10320 940 10560
rect 1180 10320 1270 10560
rect 1510 10320 1600 10560
rect 1840 10320 1930 10560
rect 2170 10320 2260 10560
rect 2500 10320 2590 10560
rect 2830 10320 2920 10560
rect 3160 10320 3250 10560
rect 3490 10320 3580 10560
rect 3820 10320 3910 10560
rect 4150 10320 4240 10560
rect 4480 10320 4570 10560
rect 4810 10320 4900 10560
rect 5140 10320 5230 10560
rect 5470 10320 5560 10560
rect 5800 10320 5890 10560
rect 6130 10320 6220 10560
rect 6460 10320 6550 10560
rect 6790 10320 6880 10560
rect 7120 10320 7260 10560
rect -4980 10230 7260 10320
rect -4980 9990 -4670 10230
rect -4430 9990 -4340 10230
rect -4100 9990 -4010 10230
rect -3770 9990 -3680 10230
rect -3440 9990 -3350 10230
rect -3110 9990 -3020 10230
rect -2780 9990 -2690 10230
rect -2450 9990 -2360 10230
rect -2120 9990 -2030 10230
rect -1790 9990 -1700 10230
rect -1460 9990 -1370 10230
rect -1130 9990 -1040 10230
rect -800 9990 -710 10230
rect -470 9990 -380 10230
rect -140 9990 -50 10230
rect 190 9990 280 10230
rect 520 9990 610 10230
rect 850 9990 940 10230
rect 1180 9990 1270 10230
rect 1510 9990 1600 10230
rect 1840 9990 1930 10230
rect 2170 9990 2260 10230
rect 2500 9990 2590 10230
rect 2830 9990 2920 10230
rect 3160 9990 3250 10230
rect 3490 9990 3580 10230
rect 3820 9990 3910 10230
rect 4150 9990 4240 10230
rect 4480 9990 4570 10230
rect 4810 9990 4900 10230
rect 5140 9990 5230 10230
rect 5470 9990 5560 10230
rect 5800 9990 5890 10230
rect 6130 9990 6220 10230
rect 6460 9990 6550 10230
rect 6790 9990 6880 10230
rect 7120 9990 7260 10230
rect -4980 9900 7260 9990
rect -4980 9660 -4670 9900
rect -4430 9660 -4340 9900
rect -4100 9660 -4010 9900
rect -3770 9660 -3680 9900
rect -3440 9660 -3350 9900
rect -3110 9660 -3020 9900
rect -2780 9660 -2690 9900
rect -2450 9660 -2360 9900
rect -2120 9660 -2030 9900
rect -1790 9660 -1700 9900
rect -1460 9660 -1370 9900
rect -1130 9660 -1040 9900
rect -800 9660 -710 9900
rect -470 9660 -380 9900
rect -140 9660 -50 9900
rect 190 9660 280 9900
rect 520 9660 610 9900
rect 850 9660 940 9900
rect 1180 9660 1270 9900
rect 1510 9660 1600 9900
rect 1840 9660 1930 9900
rect 2170 9660 2260 9900
rect 2500 9660 2590 9900
rect 2830 9660 2920 9900
rect 3160 9660 3250 9900
rect 3490 9660 3580 9900
rect 3820 9660 3910 9900
rect 4150 9660 4240 9900
rect 4480 9660 4570 9900
rect 4810 9660 4900 9900
rect 5140 9660 5230 9900
rect 5470 9660 5560 9900
rect 5800 9660 5890 9900
rect 6130 9660 6220 9900
rect 6460 9660 6550 9900
rect 6790 9660 6880 9900
rect 7120 9660 7260 9900
rect -4980 9570 7260 9660
rect -4980 9330 -4670 9570
rect -4430 9330 -4340 9570
rect -4100 9330 -4010 9570
rect -3770 9330 -3680 9570
rect -3440 9330 -3350 9570
rect -3110 9330 -3020 9570
rect -2780 9330 -2690 9570
rect -2450 9330 -2360 9570
rect -2120 9330 -2030 9570
rect -1790 9330 -1700 9570
rect -1460 9330 -1370 9570
rect -1130 9330 -1040 9570
rect -800 9330 -710 9570
rect -470 9330 -380 9570
rect -140 9330 -50 9570
rect 190 9330 280 9570
rect 520 9330 610 9570
rect 850 9330 940 9570
rect 1180 9330 1270 9570
rect 1510 9330 1600 9570
rect 1840 9330 1930 9570
rect 2170 9330 2260 9570
rect 2500 9330 2590 9570
rect 2830 9330 2920 9570
rect 3160 9330 3250 9570
rect 3490 9330 3580 9570
rect 3820 9330 3910 9570
rect 4150 9330 4240 9570
rect 4480 9330 4570 9570
rect 4810 9330 4900 9570
rect 5140 9330 5230 9570
rect 5470 9330 5560 9570
rect 5800 9330 5890 9570
rect 6130 9330 6220 9570
rect 6460 9330 6550 9570
rect 6790 9330 6880 9570
rect 7120 9330 7260 9570
rect -4980 9240 7260 9330
rect -4980 9000 -4670 9240
rect -4430 9000 -4340 9240
rect -4100 9000 -4010 9240
rect -3770 9000 -3680 9240
rect -3440 9000 -3350 9240
rect -3110 9000 -3020 9240
rect -2780 9000 -2690 9240
rect -2450 9000 -2360 9240
rect -2120 9000 -2030 9240
rect -1790 9000 -1700 9240
rect -1460 9000 -1370 9240
rect -1130 9000 -1040 9240
rect -800 9000 -710 9240
rect -470 9000 -380 9240
rect -140 9000 -50 9240
rect 190 9000 280 9240
rect 520 9000 610 9240
rect 850 9000 940 9240
rect 1180 9000 1270 9240
rect 1510 9000 1600 9240
rect 1840 9000 1930 9240
rect 2170 9000 2260 9240
rect 2500 9000 2590 9240
rect 2830 9000 2920 9240
rect 3160 9000 3250 9240
rect 3490 9000 3580 9240
rect 3820 9000 3910 9240
rect 4150 9000 4240 9240
rect 4480 9000 4570 9240
rect 4810 9000 4900 9240
rect 5140 9000 5230 9240
rect 5470 9000 5560 9240
rect 5800 9000 5890 9240
rect 6130 9000 6220 9240
rect 6460 9000 6550 9240
rect 6790 9000 6880 9240
rect 7120 9000 7260 9240
rect -4980 8870 7260 9000
rect 7640 20790 19880 21110
rect 7640 20550 7780 20790
rect 8020 20550 8110 20790
rect 8350 20550 8440 20790
rect 8680 20550 8770 20790
rect 9010 20550 9100 20790
rect 9340 20550 9430 20790
rect 9670 20550 9760 20790
rect 10000 20550 10090 20790
rect 10330 20550 10420 20790
rect 10660 20550 10750 20790
rect 10990 20550 11080 20790
rect 11320 20550 11410 20790
rect 11650 20550 11740 20790
rect 11980 20550 12070 20790
rect 12310 20550 12400 20790
rect 12640 20550 12730 20790
rect 12970 20550 13060 20790
rect 13300 20550 13390 20790
rect 13630 20550 13720 20790
rect 13960 20550 14050 20790
rect 14290 20550 14380 20790
rect 14620 20550 14710 20790
rect 14950 20550 15040 20790
rect 15280 20550 15370 20790
rect 15610 20550 15700 20790
rect 15940 20550 16030 20790
rect 16270 20550 16360 20790
rect 16600 20550 16690 20790
rect 16930 20550 17020 20790
rect 17260 20550 17350 20790
rect 17590 20550 17680 20790
rect 17920 20550 18010 20790
rect 18250 20550 18340 20790
rect 18580 20550 18670 20790
rect 18910 20550 19000 20790
rect 19240 20550 19330 20790
rect 19570 20550 19880 20790
rect 7640 20460 19880 20550
rect 7640 20220 7780 20460
rect 8020 20220 8110 20460
rect 8350 20220 8440 20460
rect 8680 20220 8770 20460
rect 9010 20220 9100 20460
rect 9340 20220 9430 20460
rect 9670 20220 9760 20460
rect 10000 20220 10090 20460
rect 10330 20220 10420 20460
rect 10660 20220 10750 20460
rect 10990 20220 11080 20460
rect 11320 20220 11410 20460
rect 11650 20220 11740 20460
rect 11980 20220 12070 20460
rect 12310 20220 12400 20460
rect 12640 20220 12730 20460
rect 12970 20220 13060 20460
rect 13300 20220 13390 20460
rect 13630 20220 13720 20460
rect 13960 20220 14050 20460
rect 14290 20220 14380 20460
rect 14620 20220 14710 20460
rect 14950 20220 15040 20460
rect 15280 20220 15370 20460
rect 15610 20220 15700 20460
rect 15940 20220 16030 20460
rect 16270 20220 16360 20460
rect 16600 20220 16690 20460
rect 16930 20220 17020 20460
rect 17260 20220 17350 20460
rect 17590 20220 17680 20460
rect 17920 20220 18010 20460
rect 18250 20220 18340 20460
rect 18580 20220 18670 20460
rect 18910 20220 19000 20460
rect 19240 20220 19330 20460
rect 19570 20220 19880 20460
rect 7640 20130 19880 20220
rect 7640 19890 7780 20130
rect 8020 19890 8110 20130
rect 8350 19890 8440 20130
rect 8680 19890 8770 20130
rect 9010 19890 9100 20130
rect 9340 19890 9430 20130
rect 9670 19890 9760 20130
rect 10000 19890 10090 20130
rect 10330 19890 10420 20130
rect 10660 19890 10750 20130
rect 10990 19890 11080 20130
rect 11320 19890 11410 20130
rect 11650 19890 11740 20130
rect 11980 19890 12070 20130
rect 12310 19890 12400 20130
rect 12640 19890 12730 20130
rect 12970 19890 13060 20130
rect 13300 19890 13390 20130
rect 13630 19890 13720 20130
rect 13960 19890 14050 20130
rect 14290 19890 14380 20130
rect 14620 19890 14710 20130
rect 14950 19890 15040 20130
rect 15280 19890 15370 20130
rect 15610 19890 15700 20130
rect 15940 19890 16030 20130
rect 16270 19890 16360 20130
rect 16600 19890 16690 20130
rect 16930 19890 17020 20130
rect 17260 19890 17350 20130
rect 17590 19890 17680 20130
rect 17920 19890 18010 20130
rect 18250 19890 18340 20130
rect 18580 19890 18670 20130
rect 18910 19890 19000 20130
rect 19240 19890 19330 20130
rect 19570 19890 19880 20130
rect 7640 19800 19880 19890
rect 7640 19560 7780 19800
rect 8020 19560 8110 19800
rect 8350 19560 8440 19800
rect 8680 19560 8770 19800
rect 9010 19560 9100 19800
rect 9340 19560 9430 19800
rect 9670 19560 9760 19800
rect 10000 19560 10090 19800
rect 10330 19560 10420 19800
rect 10660 19560 10750 19800
rect 10990 19560 11080 19800
rect 11320 19560 11410 19800
rect 11650 19560 11740 19800
rect 11980 19560 12070 19800
rect 12310 19560 12400 19800
rect 12640 19560 12730 19800
rect 12970 19560 13060 19800
rect 13300 19560 13390 19800
rect 13630 19560 13720 19800
rect 13960 19560 14050 19800
rect 14290 19560 14380 19800
rect 14620 19560 14710 19800
rect 14950 19560 15040 19800
rect 15280 19560 15370 19800
rect 15610 19560 15700 19800
rect 15940 19560 16030 19800
rect 16270 19560 16360 19800
rect 16600 19560 16690 19800
rect 16930 19560 17020 19800
rect 17260 19560 17350 19800
rect 17590 19560 17680 19800
rect 17920 19560 18010 19800
rect 18250 19560 18340 19800
rect 18580 19560 18670 19800
rect 18910 19560 19000 19800
rect 19240 19560 19330 19800
rect 19570 19560 19880 19800
rect 7640 19470 19880 19560
rect 7640 19230 7780 19470
rect 8020 19230 8110 19470
rect 8350 19230 8440 19470
rect 8680 19230 8770 19470
rect 9010 19230 9100 19470
rect 9340 19230 9430 19470
rect 9670 19230 9760 19470
rect 10000 19230 10090 19470
rect 10330 19230 10420 19470
rect 10660 19230 10750 19470
rect 10990 19230 11080 19470
rect 11320 19230 11410 19470
rect 11650 19230 11740 19470
rect 11980 19230 12070 19470
rect 12310 19230 12400 19470
rect 12640 19230 12730 19470
rect 12970 19230 13060 19470
rect 13300 19230 13390 19470
rect 13630 19230 13720 19470
rect 13960 19230 14050 19470
rect 14290 19230 14380 19470
rect 14620 19230 14710 19470
rect 14950 19230 15040 19470
rect 15280 19230 15370 19470
rect 15610 19230 15700 19470
rect 15940 19230 16030 19470
rect 16270 19230 16360 19470
rect 16600 19230 16690 19470
rect 16930 19230 17020 19470
rect 17260 19230 17350 19470
rect 17590 19230 17680 19470
rect 17920 19230 18010 19470
rect 18250 19230 18340 19470
rect 18580 19230 18670 19470
rect 18910 19230 19000 19470
rect 19240 19230 19330 19470
rect 19570 19230 19880 19470
rect 7640 19140 19880 19230
rect 7640 18900 7780 19140
rect 8020 18900 8110 19140
rect 8350 18900 8440 19140
rect 8680 18900 8770 19140
rect 9010 18900 9100 19140
rect 9340 18900 9430 19140
rect 9670 18900 9760 19140
rect 10000 18900 10090 19140
rect 10330 18900 10420 19140
rect 10660 18900 10750 19140
rect 10990 18900 11080 19140
rect 11320 18900 11410 19140
rect 11650 18900 11740 19140
rect 11980 18900 12070 19140
rect 12310 18900 12400 19140
rect 12640 18900 12730 19140
rect 12970 18900 13060 19140
rect 13300 18900 13390 19140
rect 13630 18900 13720 19140
rect 13960 18900 14050 19140
rect 14290 18900 14380 19140
rect 14620 18900 14710 19140
rect 14950 18900 15040 19140
rect 15280 18900 15370 19140
rect 15610 18900 15700 19140
rect 15940 18900 16030 19140
rect 16270 18900 16360 19140
rect 16600 18900 16690 19140
rect 16930 18900 17020 19140
rect 17260 18900 17350 19140
rect 17590 18900 17680 19140
rect 17920 18900 18010 19140
rect 18250 18900 18340 19140
rect 18580 18900 18670 19140
rect 18910 18900 19000 19140
rect 19240 18900 19330 19140
rect 19570 18900 19880 19140
rect 7640 18810 19880 18900
rect 7640 18570 7780 18810
rect 8020 18570 8110 18810
rect 8350 18570 8440 18810
rect 8680 18570 8770 18810
rect 9010 18570 9100 18810
rect 9340 18570 9430 18810
rect 9670 18570 9760 18810
rect 10000 18570 10090 18810
rect 10330 18570 10420 18810
rect 10660 18570 10750 18810
rect 10990 18570 11080 18810
rect 11320 18570 11410 18810
rect 11650 18570 11740 18810
rect 11980 18570 12070 18810
rect 12310 18570 12400 18810
rect 12640 18570 12730 18810
rect 12970 18570 13060 18810
rect 13300 18570 13390 18810
rect 13630 18570 13720 18810
rect 13960 18570 14050 18810
rect 14290 18570 14380 18810
rect 14620 18570 14710 18810
rect 14950 18570 15040 18810
rect 15280 18570 15370 18810
rect 15610 18570 15700 18810
rect 15940 18570 16030 18810
rect 16270 18570 16360 18810
rect 16600 18570 16690 18810
rect 16930 18570 17020 18810
rect 17260 18570 17350 18810
rect 17590 18570 17680 18810
rect 17920 18570 18010 18810
rect 18250 18570 18340 18810
rect 18580 18570 18670 18810
rect 18910 18570 19000 18810
rect 19240 18570 19330 18810
rect 19570 18570 19880 18810
rect 7640 18480 19880 18570
rect 7640 18240 7780 18480
rect 8020 18240 8110 18480
rect 8350 18240 8440 18480
rect 8680 18240 8770 18480
rect 9010 18240 9100 18480
rect 9340 18240 9430 18480
rect 9670 18240 9760 18480
rect 10000 18240 10090 18480
rect 10330 18240 10420 18480
rect 10660 18240 10750 18480
rect 10990 18240 11080 18480
rect 11320 18240 11410 18480
rect 11650 18240 11740 18480
rect 11980 18240 12070 18480
rect 12310 18240 12400 18480
rect 12640 18240 12730 18480
rect 12970 18240 13060 18480
rect 13300 18240 13390 18480
rect 13630 18240 13720 18480
rect 13960 18240 14050 18480
rect 14290 18240 14380 18480
rect 14620 18240 14710 18480
rect 14950 18240 15040 18480
rect 15280 18240 15370 18480
rect 15610 18240 15700 18480
rect 15940 18240 16030 18480
rect 16270 18240 16360 18480
rect 16600 18240 16690 18480
rect 16930 18240 17020 18480
rect 17260 18240 17350 18480
rect 17590 18240 17680 18480
rect 17920 18240 18010 18480
rect 18250 18240 18340 18480
rect 18580 18240 18670 18480
rect 18910 18240 19000 18480
rect 19240 18240 19330 18480
rect 19570 18240 19880 18480
rect 7640 18150 19880 18240
rect 7640 17910 7780 18150
rect 8020 17910 8110 18150
rect 8350 17910 8440 18150
rect 8680 17910 8770 18150
rect 9010 17910 9100 18150
rect 9340 17910 9430 18150
rect 9670 17910 9760 18150
rect 10000 17910 10090 18150
rect 10330 17910 10420 18150
rect 10660 17910 10750 18150
rect 10990 17910 11080 18150
rect 11320 17910 11410 18150
rect 11650 17910 11740 18150
rect 11980 17910 12070 18150
rect 12310 17910 12400 18150
rect 12640 17910 12730 18150
rect 12970 17910 13060 18150
rect 13300 17910 13390 18150
rect 13630 17910 13720 18150
rect 13960 17910 14050 18150
rect 14290 17910 14380 18150
rect 14620 17910 14710 18150
rect 14950 17910 15040 18150
rect 15280 17910 15370 18150
rect 15610 17910 15700 18150
rect 15940 17910 16030 18150
rect 16270 17910 16360 18150
rect 16600 17910 16690 18150
rect 16930 17910 17020 18150
rect 17260 17910 17350 18150
rect 17590 17910 17680 18150
rect 17920 17910 18010 18150
rect 18250 17910 18340 18150
rect 18580 17910 18670 18150
rect 18910 17910 19000 18150
rect 19240 17910 19330 18150
rect 19570 17910 19880 18150
rect 7640 17820 19880 17910
rect 7640 17580 7780 17820
rect 8020 17580 8110 17820
rect 8350 17580 8440 17820
rect 8680 17580 8770 17820
rect 9010 17580 9100 17820
rect 9340 17580 9430 17820
rect 9670 17580 9760 17820
rect 10000 17580 10090 17820
rect 10330 17580 10420 17820
rect 10660 17580 10750 17820
rect 10990 17580 11080 17820
rect 11320 17580 11410 17820
rect 11650 17580 11740 17820
rect 11980 17580 12070 17820
rect 12310 17580 12400 17820
rect 12640 17580 12730 17820
rect 12970 17580 13060 17820
rect 13300 17580 13390 17820
rect 13630 17580 13720 17820
rect 13960 17580 14050 17820
rect 14290 17580 14380 17820
rect 14620 17580 14710 17820
rect 14950 17580 15040 17820
rect 15280 17580 15370 17820
rect 15610 17580 15700 17820
rect 15940 17580 16030 17820
rect 16270 17580 16360 17820
rect 16600 17580 16690 17820
rect 16930 17580 17020 17820
rect 17260 17580 17350 17820
rect 17590 17580 17680 17820
rect 17920 17580 18010 17820
rect 18250 17580 18340 17820
rect 18580 17580 18670 17820
rect 18910 17580 19000 17820
rect 19240 17580 19330 17820
rect 19570 17580 19880 17820
rect 7640 17490 19880 17580
rect 7640 17250 7780 17490
rect 8020 17250 8110 17490
rect 8350 17250 8440 17490
rect 8680 17250 8770 17490
rect 9010 17250 9100 17490
rect 9340 17250 9430 17490
rect 9670 17250 9760 17490
rect 10000 17250 10090 17490
rect 10330 17250 10420 17490
rect 10660 17250 10750 17490
rect 10990 17250 11080 17490
rect 11320 17250 11410 17490
rect 11650 17250 11740 17490
rect 11980 17250 12070 17490
rect 12310 17250 12400 17490
rect 12640 17250 12730 17490
rect 12970 17250 13060 17490
rect 13300 17250 13390 17490
rect 13630 17250 13720 17490
rect 13960 17250 14050 17490
rect 14290 17250 14380 17490
rect 14620 17250 14710 17490
rect 14950 17250 15040 17490
rect 15280 17250 15370 17490
rect 15610 17250 15700 17490
rect 15940 17250 16030 17490
rect 16270 17250 16360 17490
rect 16600 17250 16690 17490
rect 16930 17250 17020 17490
rect 17260 17250 17350 17490
rect 17590 17250 17680 17490
rect 17920 17250 18010 17490
rect 18250 17250 18340 17490
rect 18580 17250 18670 17490
rect 18910 17250 19000 17490
rect 19240 17250 19330 17490
rect 19570 17250 19880 17490
rect 7640 17160 19880 17250
rect 7640 16920 7780 17160
rect 8020 16920 8110 17160
rect 8350 16920 8440 17160
rect 8680 16920 8770 17160
rect 9010 16920 9100 17160
rect 9340 16920 9430 17160
rect 9670 16920 9760 17160
rect 10000 16920 10090 17160
rect 10330 16920 10420 17160
rect 10660 16920 10750 17160
rect 10990 16920 11080 17160
rect 11320 16920 11410 17160
rect 11650 16920 11740 17160
rect 11980 16920 12070 17160
rect 12310 16920 12400 17160
rect 12640 16920 12730 17160
rect 12970 16920 13060 17160
rect 13300 16920 13390 17160
rect 13630 16920 13720 17160
rect 13960 16920 14050 17160
rect 14290 16920 14380 17160
rect 14620 16920 14710 17160
rect 14950 16920 15040 17160
rect 15280 16920 15370 17160
rect 15610 16920 15700 17160
rect 15940 16920 16030 17160
rect 16270 16920 16360 17160
rect 16600 16920 16690 17160
rect 16930 16920 17020 17160
rect 17260 16920 17350 17160
rect 17590 16920 17680 17160
rect 17920 16920 18010 17160
rect 18250 16920 18340 17160
rect 18580 16920 18670 17160
rect 18910 16920 19000 17160
rect 19240 16920 19330 17160
rect 19570 16920 19880 17160
rect 7640 16830 19880 16920
rect 7640 16590 7780 16830
rect 8020 16590 8110 16830
rect 8350 16590 8440 16830
rect 8680 16590 8770 16830
rect 9010 16590 9100 16830
rect 9340 16590 9430 16830
rect 9670 16590 9760 16830
rect 10000 16590 10090 16830
rect 10330 16590 10420 16830
rect 10660 16590 10750 16830
rect 10990 16590 11080 16830
rect 11320 16590 11410 16830
rect 11650 16590 11740 16830
rect 11980 16590 12070 16830
rect 12310 16590 12400 16830
rect 12640 16590 12730 16830
rect 12970 16590 13060 16830
rect 13300 16590 13390 16830
rect 13630 16590 13720 16830
rect 13960 16590 14050 16830
rect 14290 16590 14380 16830
rect 14620 16590 14710 16830
rect 14950 16590 15040 16830
rect 15280 16590 15370 16830
rect 15610 16590 15700 16830
rect 15940 16590 16030 16830
rect 16270 16590 16360 16830
rect 16600 16590 16690 16830
rect 16930 16590 17020 16830
rect 17260 16590 17350 16830
rect 17590 16590 17680 16830
rect 17920 16590 18010 16830
rect 18250 16590 18340 16830
rect 18580 16590 18670 16830
rect 18910 16590 19000 16830
rect 19240 16590 19330 16830
rect 19570 16590 19880 16830
rect 7640 16500 19880 16590
rect 7640 16260 7780 16500
rect 8020 16260 8110 16500
rect 8350 16260 8440 16500
rect 8680 16260 8770 16500
rect 9010 16260 9100 16500
rect 9340 16260 9430 16500
rect 9670 16260 9760 16500
rect 10000 16260 10090 16500
rect 10330 16260 10420 16500
rect 10660 16260 10750 16500
rect 10990 16260 11080 16500
rect 11320 16260 11410 16500
rect 11650 16260 11740 16500
rect 11980 16260 12070 16500
rect 12310 16260 12400 16500
rect 12640 16260 12730 16500
rect 12970 16260 13060 16500
rect 13300 16260 13390 16500
rect 13630 16260 13720 16500
rect 13960 16260 14050 16500
rect 14290 16260 14380 16500
rect 14620 16260 14710 16500
rect 14950 16260 15040 16500
rect 15280 16260 15370 16500
rect 15610 16260 15700 16500
rect 15940 16260 16030 16500
rect 16270 16260 16360 16500
rect 16600 16260 16690 16500
rect 16930 16260 17020 16500
rect 17260 16260 17350 16500
rect 17590 16260 17680 16500
rect 17920 16260 18010 16500
rect 18250 16260 18340 16500
rect 18580 16260 18670 16500
rect 18910 16260 19000 16500
rect 19240 16260 19330 16500
rect 19570 16260 19880 16500
rect 7640 16170 19880 16260
rect 7640 15930 7780 16170
rect 8020 15930 8110 16170
rect 8350 15930 8440 16170
rect 8680 15930 8770 16170
rect 9010 15930 9100 16170
rect 9340 15930 9430 16170
rect 9670 15930 9760 16170
rect 10000 15930 10090 16170
rect 10330 15930 10420 16170
rect 10660 15930 10750 16170
rect 10990 15930 11080 16170
rect 11320 15930 11410 16170
rect 11650 15930 11740 16170
rect 11980 15930 12070 16170
rect 12310 15930 12400 16170
rect 12640 15930 12730 16170
rect 12970 15930 13060 16170
rect 13300 15930 13390 16170
rect 13630 15930 13720 16170
rect 13960 15930 14050 16170
rect 14290 15930 14380 16170
rect 14620 15930 14710 16170
rect 14950 15930 15040 16170
rect 15280 15930 15370 16170
rect 15610 15930 15700 16170
rect 15940 15930 16030 16170
rect 16270 15930 16360 16170
rect 16600 15930 16690 16170
rect 16930 15930 17020 16170
rect 17260 15930 17350 16170
rect 17590 15930 17680 16170
rect 17920 15930 18010 16170
rect 18250 15930 18340 16170
rect 18580 15930 18670 16170
rect 18910 15930 19000 16170
rect 19240 15930 19330 16170
rect 19570 15930 19880 16170
rect 7640 15840 19880 15930
rect 7640 15600 7780 15840
rect 8020 15600 8110 15840
rect 8350 15600 8440 15840
rect 8680 15600 8770 15840
rect 9010 15600 9100 15840
rect 9340 15600 9430 15840
rect 9670 15600 9760 15840
rect 10000 15600 10090 15840
rect 10330 15600 10420 15840
rect 10660 15600 10750 15840
rect 10990 15600 11080 15840
rect 11320 15600 11410 15840
rect 11650 15600 11740 15840
rect 11980 15600 12070 15840
rect 12310 15600 12400 15840
rect 12640 15600 12730 15840
rect 12970 15600 13060 15840
rect 13300 15600 13390 15840
rect 13630 15600 13720 15840
rect 13960 15600 14050 15840
rect 14290 15600 14380 15840
rect 14620 15600 14710 15840
rect 14950 15600 15040 15840
rect 15280 15600 15370 15840
rect 15610 15600 15700 15840
rect 15940 15600 16030 15840
rect 16270 15600 16360 15840
rect 16600 15600 16690 15840
rect 16930 15600 17020 15840
rect 17260 15600 17350 15840
rect 17590 15600 17680 15840
rect 17920 15600 18010 15840
rect 18250 15600 18340 15840
rect 18580 15600 18670 15840
rect 18910 15600 19000 15840
rect 19240 15600 19330 15840
rect 19570 15600 19880 15840
rect 7640 15510 19880 15600
rect 7640 15270 7780 15510
rect 8020 15270 8110 15510
rect 8350 15270 8440 15510
rect 8680 15270 8770 15510
rect 9010 15270 9100 15510
rect 9340 15270 9430 15510
rect 9670 15270 9760 15510
rect 10000 15270 10090 15510
rect 10330 15270 10420 15510
rect 10660 15270 10750 15510
rect 10990 15270 11080 15510
rect 11320 15270 11410 15510
rect 11650 15270 11740 15510
rect 11980 15270 12070 15510
rect 12310 15270 12400 15510
rect 12640 15270 12730 15510
rect 12970 15270 13060 15510
rect 13300 15270 13390 15510
rect 13630 15270 13720 15510
rect 13960 15270 14050 15510
rect 14290 15270 14380 15510
rect 14620 15270 14710 15510
rect 14950 15270 15040 15510
rect 15280 15270 15370 15510
rect 15610 15270 15700 15510
rect 15940 15270 16030 15510
rect 16270 15270 16360 15510
rect 16600 15270 16690 15510
rect 16930 15270 17020 15510
rect 17260 15270 17350 15510
rect 17590 15270 17680 15510
rect 17920 15270 18010 15510
rect 18250 15270 18340 15510
rect 18580 15270 18670 15510
rect 18910 15270 19000 15510
rect 19240 15270 19330 15510
rect 19570 15270 19880 15510
rect 7640 15180 19880 15270
rect 7640 14940 7780 15180
rect 8020 14940 8110 15180
rect 8350 14940 8440 15180
rect 8680 14940 8770 15180
rect 9010 14940 9100 15180
rect 9340 14940 9430 15180
rect 9670 14940 9760 15180
rect 10000 14940 10090 15180
rect 10330 14940 10420 15180
rect 10660 14940 10750 15180
rect 10990 14940 11080 15180
rect 11320 14940 11410 15180
rect 11650 14940 11740 15180
rect 11980 14940 12070 15180
rect 12310 14940 12400 15180
rect 12640 14940 12730 15180
rect 12970 14940 13060 15180
rect 13300 14940 13390 15180
rect 13630 14940 13720 15180
rect 13960 14940 14050 15180
rect 14290 14940 14380 15180
rect 14620 14940 14710 15180
rect 14950 14940 15040 15180
rect 15280 14940 15370 15180
rect 15610 14940 15700 15180
rect 15940 14940 16030 15180
rect 16270 14940 16360 15180
rect 16600 14940 16690 15180
rect 16930 14940 17020 15180
rect 17260 14940 17350 15180
rect 17590 14940 17680 15180
rect 17920 14940 18010 15180
rect 18250 14940 18340 15180
rect 18580 14940 18670 15180
rect 18910 14940 19000 15180
rect 19240 14940 19330 15180
rect 19570 14940 19880 15180
rect 7640 14850 19880 14940
rect 7640 14610 7780 14850
rect 8020 14610 8110 14850
rect 8350 14610 8440 14850
rect 8680 14610 8770 14850
rect 9010 14610 9100 14850
rect 9340 14610 9430 14850
rect 9670 14610 9760 14850
rect 10000 14610 10090 14850
rect 10330 14610 10420 14850
rect 10660 14610 10750 14850
rect 10990 14610 11080 14850
rect 11320 14610 11410 14850
rect 11650 14610 11740 14850
rect 11980 14610 12070 14850
rect 12310 14610 12400 14850
rect 12640 14610 12730 14850
rect 12970 14610 13060 14850
rect 13300 14610 13390 14850
rect 13630 14610 13720 14850
rect 13960 14610 14050 14850
rect 14290 14610 14380 14850
rect 14620 14610 14710 14850
rect 14950 14610 15040 14850
rect 15280 14610 15370 14850
rect 15610 14610 15700 14850
rect 15940 14610 16030 14850
rect 16270 14610 16360 14850
rect 16600 14610 16690 14850
rect 16930 14610 17020 14850
rect 17260 14610 17350 14850
rect 17590 14610 17680 14850
rect 17920 14610 18010 14850
rect 18250 14610 18340 14850
rect 18580 14610 18670 14850
rect 18910 14610 19000 14850
rect 19240 14610 19330 14850
rect 19570 14610 19880 14850
rect 7640 14520 19880 14610
rect 7640 14280 7780 14520
rect 8020 14280 8110 14520
rect 8350 14280 8440 14520
rect 8680 14280 8770 14520
rect 9010 14280 9100 14520
rect 9340 14280 9430 14520
rect 9670 14280 9760 14520
rect 10000 14280 10090 14520
rect 10330 14280 10420 14520
rect 10660 14280 10750 14520
rect 10990 14280 11080 14520
rect 11320 14280 11410 14520
rect 11650 14280 11740 14520
rect 11980 14280 12070 14520
rect 12310 14280 12400 14520
rect 12640 14280 12730 14520
rect 12970 14280 13060 14520
rect 13300 14280 13390 14520
rect 13630 14280 13720 14520
rect 13960 14280 14050 14520
rect 14290 14280 14380 14520
rect 14620 14280 14710 14520
rect 14950 14280 15040 14520
rect 15280 14280 15370 14520
rect 15610 14280 15700 14520
rect 15940 14280 16030 14520
rect 16270 14280 16360 14520
rect 16600 14280 16690 14520
rect 16930 14280 17020 14520
rect 17260 14280 17350 14520
rect 17590 14280 17680 14520
rect 17920 14280 18010 14520
rect 18250 14280 18340 14520
rect 18580 14280 18670 14520
rect 18910 14280 19000 14520
rect 19240 14280 19330 14520
rect 19570 14280 19880 14520
rect 7640 14190 19880 14280
rect 7640 13950 7780 14190
rect 8020 13950 8110 14190
rect 8350 13950 8440 14190
rect 8680 13950 8770 14190
rect 9010 13950 9100 14190
rect 9340 13950 9430 14190
rect 9670 13950 9760 14190
rect 10000 13950 10090 14190
rect 10330 13950 10420 14190
rect 10660 13950 10750 14190
rect 10990 13950 11080 14190
rect 11320 13950 11410 14190
rect 11650 13950 11740 14190
rect 11980 13950 12070 14190
rect 12310 13950 12400 14190
rect 12640 13950 12730 14190
rect 12970 13950 13060 14190
rect 13300 13950 13390 14190
rect 13630 13950 13720 14190
rect 13960 13950 14050 14190
rect 14290 13950 14380 14190
rect 14620 13950 14710 14190
rect 14950 13950 15040 14190
rect 15280 13950 15370 14190
rect 15610 13950 15700 14190
rect 15940 13950 16030 14190
rect 16270 13950 16360 14190
rect 16600 13950 16690 14190
rect 16930 13950 17020 14190
rect 17260 13950 17350 14190
rect 17590 13950 17680 14190
rect 17920 13950 18010 14190
rect 18250 13950 18340 14190
rect 18580 13950 18670 14190
rect 18910 13950 19000 14190
rect 19240 13950 19330 14190
rect 19570 13950 19880 14190
rect 7640 13860 19880 13950
rect 7640 13620 7780 13860
rect 8020 13620 8110 13860
rect 8350 13620 8440 13860
rect 8680 13620 8770 13860
rect 9010 13620 9100 13860
rect 9340 13620 9430 13860
rect 9670 13620 9760 13860
rect 10000 13620 10090 13860
rect 10330 13620 10420 13860
rect 10660 13620 10750 13860
rect 10990 13620 11080 13860
rect 11320 13620 11410 13860
rect 11650 13620 11740 13860
rect 11980 13620 12070 13860
rect 12310 13620 12400 13860
rect 12640 13620 12730 13860
rect 12970 13620 13060 13860
rect 13300 13620 13390 13860
rect 13630 13620 13720 13860
rect 13960 13620 14050 13860
rect 14290 13620 14380 13860
rect 14620 13620 14710 13860
rect 14950 13620 15040 13860
rect 15280 13620 15370 13860
rect 15610 13620 15700 13860
rect 15940 13620 16030 13860
rect 16270 13620 16360 13860
rect 16600 13620 16690 13860
rect 16930 13620 17020 13860
rect 17260 13620 17350 13860
rect 17590 13620 17680 13860
rect 17920 13620 18010 13860
rect 18250 13620 18340 13860
rect 18580 13620 18670 13860
rect 18910 13620 19000 13860
rect 19240 13620 19330 13860
rect 19570 13620 19880 13860
rect 7640 13530 19880 13620
rect 7640 13290 7780 13530
rect 8020 13290 8110 13530
rect 8350 13290 8440 13530
rect 8680 13290 8770 13530
rect 9010 13290 9100 13530
rect 9340 13290 9430 13530
rect 9670 13290 9760 13530
rect 10000 13290 10090 13530
rect 10330 13290 10420 13530
rect 10660 13290 10750 13530
rect 10990 13290 11080 13530
rect 11320 13290 11410 13530
rect 11650 13290 11740 13530
rect 11980 13290 12070 13530
rect 12310 13290 12400 13530
rect 12640 13290 12730 13530
rect 12970 13290 13060 13530
rect 13300 13290 13390 13530
rect 13630 13290 13720 13530
rect 13960 13290 14050 13530
rect 14290 13290 14380 13530
rect 14620 13290 14710 13530
rect 14950 13290 15040 13530
rect 15280 13290 15370 13530
rect 15610 13290 15700 13530
rect 15940 13290 16030 13530
rect 16270 13290 16360 13530
rect 16600 13290 16690 13530
rect 16930 13290 17020 13530
rect 17260 13290 17350 13530
rect 17590 13290 17680 13530
rect 17920 13290 18010 13530
rect 18250 13290 18340 13530
rect 18580 13290 18670 13530
rect 18910 13290 19000 13530
rect 19240 13290 19330 13530
rect 19570 13290 19880 13530
rect 7640 13200 19880 13290
rect 7640 12960 7780 13200
rect 8020 12960 8110 13200
rect 8350 12960 8440 13200
rect 8680 12960 8770 13200
rect 9010 12960 9100 13200
rect 9340 12960 9430 13200
rect 9670 12960 9760 13200
rect 10000 12960 10090 13200
rect 10330 12960 10420 13200
rect 10660 12960 10750 13200
rect 10990 12960 11080 13200
rect 11320 12960 11410 13200
rect 11650 12960 11740 13200
rect 11980 12960 12070 13200
rect 12310 12960 12400 13200
rect 12640 12960 12730 13200
rect 12970 12960 13060 13200
rect 13300 12960 13390 13200
rect 13630 12960 13720 13200
rect 13960 12960 14050 13200
rect 14290 12960 14380 13200
rect 14620 12960 14710 13200
rect 14950 12960 15040 13200
rect 15280 12960 15370 13200
rect 15610 12960 15700 13200
rect 15940 12960 16030 13200
rect 16270 12960 16360 13200
rect 16600 12960 16690 13200
rect 16930 12960 17020 13200
rect 17260 12960 17350 13200
rect 17590 12960 17680 13200
rect 17920 12960 18010 13200
rect 18250 12960 18340 13200
rect 18580 12960 18670 13200
rect 18910 12960 19000 13200
rect 19240 12960 19330 13200
rect 19570 12960 19880 13200
rect 7640 12870 19880 12960
rect 7640 12630 7780 12870
rect 8020 12630 8110 12870
rect 8350 12630 8440 12870
rect 8680 12630 8770 12870
rect 9010 12630 9100 12870
rect 9340 12630 9430 12870
rect 9670 12630 9760 12870
rect 10000 12630 10090 12870
rect 10330 12630 10420 12870
rect 10660 12630 10750 12870
rect 10990 12630 11080 12870
rect 11320 12630 11410 12870
rect 11650 12630 11740 12870
rect 11980 12630 12070 12870
rect 12310 12630 12400 12870
rect 12640 12630 12730 12870
rect 12970 12630 13060 12870
rect 13300 12630 13390 12870
rect 13630 12630 13720 12870
rect 13960 12630 14050 12870
rect 14290 12630 14380 12870
rect 14620 12630 14710 12870
rect 14950 12630 15040 12870
rect 15280 12630 15370 12870
rect 15610 12630 15700 12870
rect 15940 12630 16030 12870
rect 16270 12630 16360 12870
rect 16600 12630 16690 12870
rect 16930 12630 17020 12870
rect 17260 12630 17350 12870
rect 17590 12630 17680 12870
rect 17920 12630 18010 12870
rect 18250 12630 18340 12870
rect 18580 12630 18670 12870
rect 18910 12630 19000 12870
rect 19240 12630 19330 12870
rect 19570 12630 19880 12870
rect 7640 12540 19880 12630
rect 7640 12300 7780 12540
rect 8020 12300 8110 12540
rect 8350 12300 8440 12540
rect 8680 12300 8770 12540
rect 9010 12300 9100 12540
rect 9340 12300 9430 12540
rect 9670 12300 9760 12540
rect 10000 12300 10090 12540
rect 10330 12300 10420 12540
rect 10660 12300 10750 12540
rect 10990 12300 11080 12540
rect 11320 12300 11410 12540
rect 11650 12300 11740 12540
rect 11980 12300 12070 12540
rect 12310 12300 12400 12540
rect 12640 12300 12730 12540
rect 12970 12300 13060 12540
rect 13300 12300 13390 12540
rect 13630 12300 13720 12540
rect 13960 12300 14050 12540
rect 14290 12300 14380 12540
rect 14620 12300 14710 12540
rect 14950 12300 15040 12540
rect 15280 12300 15370 12540
rect 15610 12300 15700 12540
rect 15940 12300 16030 12540
rect 16270 12300 16360 12540
rect 16600 12300 16690 12540
rect 16930 12300 17020 12540
rect 17260 12300 17350 12540
rect 17590 12300 17680 12540
rect 17920 12300 18010 12540
rect 18250 12300 18340 12540
rect 18580 12300 18670 12540
rect 18910 12300 19000 12540
rect 19240 12300 19330 12540
rect 19570 12300 19880 12540
rect 7640 12210 19880 12300
rect 7640 11970 7780 12210
rect 8020 11970 8110 12210
rect 8350 11970 8440 12210
rect 8680 11970 8770 12210
rect 9010 11970 9100 12210
rect 9340 11970 9430 12210
rect 9670 11970 9760 12210
rect 10000 11970 10090 12210
rect 10330 11970 10420 12210
rect 10660 11970 10750 12210
rect 10990 11970 11080 12210
rect 11320 11970 11410 12210
rect 11650 11970 11740 12210
rect 11980 11970 12070 12210
rect 12310 11970 12400 12210
rect 12640 11970 12730 12210
rect 12970 11970 13060 12210
rect 13300 11970 13390 12210
rect 13630 11970 13720 12210
rect 13960 11970 14050 12210
rect 14290 11970 14380 12210
rect 14620 11970 14710 12210
rect 14950 11970 15040 12210
rect 15280 11970 15370 12210
rect 15610 11970 15700 12210
rect 15940 11970 16030 12210
rect 16270 11970 16360 12210
rect 16600 11970 16690 12210
rect 16930 11970 17020 12210
rect 17260 11970 17350 12210
rect 17590 11970 17680 12210
rect 17920 11970 18010 12210
rect 18250 11970 18340 12210
rect 18580 11970 18670 12210
rect 18910 11970 19000 12210
rect 19240 11970 19330 12210
rect 19570 11970 19880 12210
rect 7640 11880 19880 11970
rect 7640 11640 7780 11880
rect 8020 11640 8110 11880
rect 8350 11640 8440 11880
rect 8680 11640 8770 11880
rect 9010 11640 9100 11880
rect 9340 11640 9430 11880
rect 9670 11640 9760 11880
rect 10000 11640 10090 11880
rect 10330 11640 10420 11880
rect 10660 11640 10750 11880
rect 10990 11640 11080 11880
rect 11320 11640 11410 11880
rect 11650 11640 11740 11880
rect 11980 11640 12070 11880
rect 12310 11640 12400 11880
rect 12640 11640 12730 11880
rect 12970 11640 13060 11880
rect 13300 11640 13390 11880
rect 13630 11640 13720 11880
rect 13960 11640 14050 11880
rect 14290 11640 14380 11880
rect 14620 11640 14710 11880
rect 14950 11640 15040 11880
rect 15280 11640 15370 11880
rect 15610 11640 15700 11880
rect 15940 11640 16030 11880
rect 16270 11640 16360 11880
rect 16600 11640 16690 11880
rect 16930 11640 17020 11880
rect 17260 11640 17350 11880
rect 17590 11640 17680 11880
rect 17920 11640 18010 11880
rect 18250 11640 18340 11880
rect 18580 11640 18670 11880
rect 18910 11640 19000 11880
rect 19240 11640 19330 11880
rect 19570 11640 19880 11880
rect 7640 11550 19880 11640
rect 7640 11310 7780 11550
rect 8020 11310 8110 11550
rect 8350 11310 8440 11550
rect 8680 11310 8770 11550
rect 9010 11310 9100 11550
rect 9340 11310 9430 11550
rect 9670 11310 9760 11550
rect 10000 11310 10090 11550
rect 10330 11310 10420 11550
rect 10660 11310 10750 11550
rect 10990 11310 11080 11550
rect 11320 11310 11410 11550
rect 11650 11310 11740 11550
rect 11980 11310 12070 11550
rect 12310 11310 12400 11550
rect 12640 11310 12730 11550
rect 12970 11310 13060 11550
rect 13300 11310 13390 11550
rect 13630 11310 13720 11550
rect 13960 11310 14050 11550
rect 14290 11310 14380 11550
rect 14620 11310 14710 11550
rect 14950 11310 15040 11550
rect 15280 11310 15370 11550
rect 15610 11310 15700 11550
rect 15940 11310 16030 11550
rect 16270 11310 16360 11550
rect 16600 11310 16690 11550
rect 16930 11310 17020 11550
rect 17260 11310 17350 11550
rect 17590 11310 17680 11550
rect 17920 11310 18010 11550
rect 18250 11310 18340 11550
rect 18580 11310 18670 11550
rect 18910 11310 19000 11550
rect 19240 11310 19330 11550
rect 19570 11310 19880 11550
rect 7640 11220 19880 11310
rect 7640 10980 7780 11220
rect 8020 10980 8110 11220
rect 8350 10980 8440 11220
rect 8680 10980 8770 11220
rect 9010 10980 9100 11220
rect 9340 10980 9430 11220
rect 9670 10980 9760 11220
rect 10000 10980 10090 11220
rect 10330 10980 10420 11220
rect 10660 10980 10750 11220
rect 10990 10980 11080 11220
rect 11320 10980 11410 11220
rect 11650 10980 11740 11220
rect 11980 10980 12070 11220
rect 12310 10980 12400 11220
rect 12640 10980 12730 11220
rect 12970 10980 13060 11220
rect 13300 10980 13390 11220
rect 13630 10980 13720 11220
rect 13960 10980 14050 11220
rect 14290 10980 14380 11220
rect 14620 10980 14710 11220
rect 14950 10980 15040 11220
rect 15280 10980 15370 11220
rect 15610 10980 15700 11220
rect 15940 10980 16030 11220
rect 16270 10980 16360 11220
rect 16600 10980 16690 11220
rect 16930 10980 17020 11220
rect 17260 10980 17350 11220
rect 17590 10980 17680 11220
rect 17920 10980 18010 11220
rect 18250 10980 18340 11220
rect 18580 10980 18670 11220
rect 18910 10980 19000 11220
rect 19240 10980 19330 11220
rect 19570 10980 19880 11220
rect 7640 10890 19880 10980
rect 7640 10650 7780 10890
rect 8020 10650 8110 10890
rect 8350 10650 8440 10890
rect 8680 10650 8770 10890
rect 9010 10650 9100 10890
rect 9340 10650 9430 10890
rect 9670 10650 9760 10890
rect 10000 10650 10090 10890
rect 10330 10650 10420 10890
rect 10660 10650 10750 10890
rect 10990 10650 11080 10890
rect 11320 10650 11410 10890
rect 11650 10650 11740 10890
rect 11980 10650 12070 10890
rect 12310 10650 12400 10890
rect 12640 10650 12730 10890
rect 12970 10650 13060 10890
rect 13300 10650 13390 10890
rect 13630 10650 13720 10890
rect 13960 10650 14050 10890
rect 14290 10650 14380 10890
rect 14620 10650 14710 10890
rect 14950 10650 15040 10890
rect 15280 10650 15370 10890
rect 15610 10650 15700 10890
rect 15940 10650 16030 10890
rect 16270 10650 16360 10890
rect 16600 10650 16690 10890
rect 16930 10650 17020 10890
rect 17260 10650 17350 10890
rect 17590 10650 17680 10890
rect 17920 10650 18010 10890
rect 18250 10650 18340 10890
rect 18580 10650 18670 10890
rect 18910 10650 19000 10890
rect 19240 10650 19330 10890
rect 19570 10650 19880 10890
rect 7640 10560 19880 10650
rect 7640 10320 7780 10560
rect 8020 10320 8110 10560
rect 8350 10320 8440 10560
rect 8680 10320 8770 10560
rect 9010 10320 9100 10560
rect 9340 10320 9430 10560
rect 9670 10320 9760 10560
rect 10000 10320 10090 10560
rect 10330 10320 10420 10560
rect 10660 10320 10750 10560
rect 10990 10320 11080 10560
rect 11320 10320 11410 10560
rect 11650 10320 11740 10560
rect 11980 10320 12070 10560
rect 12310 10320 12400 10560
rect 12640 10320 12730 10560
rect 12970 10320 13060 10560
rect 13300 10320 13390 10560
rect 13630 10320 13720 10560
rect 13960 10320 14050 10560
rect 14290 10320 14380 10560
rect 14620 10320 14710 10560
rect 14950 10320 15040 10560
rect 15280 10320 15370 10560
rect 15610 10320 15700 10560
rect 15940 10320 16030 10560
rect 16270 10320 16360 10560
rect 16600 10320 16690 10560
rect 16930 10320 17020 10560
rect 17260 10320 17350 10560
rect 17590 10320 17680 10560
rect 17920 10320 18010 10560
rect 18250 10320 18340 10560
rect 18580 10320 18670 10560
rect 18910 10320 19000 10560
rect 19240 10320 19330 10560
rect 19570 10320 19880 10560
rect 7640 10230 19880 10320
rect 7640 9990 7780 10230
rect 8020 9990 8110 10230
rect 8350 9990 8440 10230
rect 8680 9990 8770 10230
rect 9010 9990 9100 10230
rect 9340 9990 9430 10230
rect 9670 9990 9760 10230
rect 10000 9990 10090 10230
rect 10330 9990 10420 10230
rect 10660 9990 10750 10230
rect 10990 9990 11080 10230
rect 11320 9990 11410 10230
rect 11650 9990 11740 10230
rect 11980 9990 12070 10230
rect 12310 9990 12400 10230
rect 12640 9990 12730 10230
rect 12970 9990 13060 10230
rect 13300 9990 13390 10230
rect 13630 9990 13720 10230
rect 13960 9990 14050 10230
rect 14290 9990 14380 10230
rect 14620 9990 14710 10230
rect 14950 9990 15040 10230
rect 15280 9990 15370 10230
rect 15610 9990 15700 10230
rect 15940 9990 16030 10230
rect 16270 9990 16360 10230
rect 16600 9990 16690 10230
rect 16930 9990 17020 10230
rect 17260 9990 17350 10230
rect 17590 9990 17680 10230
rect 17920 9990 18010 10230
rect 18250 9990 18340 10230
rect 18580 9990 18670 10230
rect 18910 9990 19000 10230
rect 19240 9990 19330 10230
rect 19570 9990 19880 10230
rect 7640 9900 19880 9990
rect 7640 9660 7780 9900
rect 8020 9660 8110 9900
rect 8350 9660 8440 9900
rect 8680 9660 8770 9900
rect 9010 9660 9100 9900
rect 9340 9660 9430 9900
rect 9670 9660 9760 9900
rect 10000 9660 10090 9900
rect 10330 9660 10420 9900
rect 10660 9660 10750 9900
rect 10990 9660 11080 9900
rect 11320 9660 11410 9900
rect 11650 9660 11740 9900
rect 11980 9660 12070 9900
rect 12310 9660 12400 9900
rect 12640 9660 12730 9900
rect 12970 9660 13060 9900
rect 13300 9660 13390 9900
rect 13630 9660 13720 9900
rect 13960 9660 14050 9900
rect 14290 9660 14380 9900
rect 14620 9660 14710 9900
rect 14950 9660 15040 9900
rect 15280 9660 15370 9900
rect 15610 9660 15700 9900
rect 15940 9660 16030 9900
rect 16270 9660 16360 9900
rect 16600 9660 16690 9900
rect 16930 9660 17020 9900
rect 17260 9660 17350 9900
rect 17590 9660 17680 9900
rect 17920 9660 18010 9900
rect 18250 9660 18340 9900
rect 18580 9660 18670 9900
rect 18910 9660 19000 9900
rect 19240 9660 19330 9900
rect 19570 9660 19880 9900
rect 7640 9570 19880 9660
rect 7640 9330 7780 9570
rect 8020 9330 8110 9570
rect 8350 9330 8440 9570
rect 8680 9330 8770 9570
rect 9010 9330 9100 9570
rect 9340 9330 9430 9570
rect 9670 9330 9760 9570
rect 10000 9330 10090 9570
rect 10330 9330 10420 9570
rect 10660 9330 10750 9570
rect 10990 9330 11080 9570
rect 11320 9330 11410 9570
rect 11650 9330 11740 9570
rect 11980 9330 12070 9570
rect 12310 9330 12400 9570
rect 12640 9330 12730 9570
rect 12970 9330 13060 9570
rect 13300 9330 13390 9570
rect 13630 9330 13720 9570
rect 13960 9330 14050 9570
rect 14290 9330 14380 9570
rect 14620 9330 14710 9570
rect 14950 9330 15040 9570
rect 15280 9330 15370 9570
rect 15610 9330 15700 9570
rect 15940 9330 16030 9570
rect 16270 9330 16360 9570
rect 16600 9330 16690 9570
rect 16930 9330 17020 9570
rect 17260 9330 17350 9570
rect 17590 9330 17680 9570
rect 17920 9330 18010 9570
rect 18250 9330 18340 9570
rect 18580 9330 18670 9570
rect 18910 9330 19000 9570
rect 19240 9330 19330 9570
rect 19570 9330 19880 9570
rect 7640 9240 19880 9330
rect 7640 9000 7780 9240
rect 8020 9000 8110 9240
rect 8350 9000 8440 9240
rect 8680 9000 8770 9240
rect 9010 9000 9100 9240
rect 9340 9000 9430 9240
rect 9670 9000 9760 9240
rect 10000 9000 10090 9240
rect 10330 9000 10420 9240
rect 10660 9000 10750 9240
rect 10990 9000 11080 9240
rect 11320 9000 11410 9240
rect 11650 9000 11740 9240
rect 11980 9000 12070 9240
rect 12310 9000 12400 9240
rect 12640 9000 12730 9240
rect 12970 9000 13060 9240
rect 13300 9000 13390 9240
rect 13630 9000 13720 9240
rect 13960 9000 14050 9240
rect 14290 9000 14380 9240
rect 14620 9000 14710 9240
rect 14950 9000 15040 9240
rect 15280 9000 15370 9240
rect 15610 9000 15700 9240
rect 15940 9000 16030 9240
rect 16270 9000 16360 9240
rect 16600 9000 16690 9240
rect 16930 9000 17020 9240
rect 17260 9000 17350 9240
rect 17590 9000 17680 9240
rect 17920 9000 18010 9240
rect 18250 9000 18340 9240
rect 18580 9000 18670 9240
rect 18910 9000 19000 9240
rect 19240 9000 19330 9240
rect 19570 9000 19880 9240
rect 7640 8870 19880 9000
rect 28730 7830 35430 7880
rect 28730 7590 28780 7830
rect 29020 7590 29110 7830
rect 29350 7590 29440 7830
rect 29680 7590 29770 7830
rect 30010 7590 30100 7830
rect 30340 7590 30430 7830
rect 30670 7590 30760 7830
rect 31000 7590 31090 7830
rect 31330 7590 31420 7830
rect 31660 7590 31750 7830
rect 31990 7590 32080 7830
rect 32320 7590 32410 7830
rect 32650 7590 32740 7830
rect 32980 7590 33070 7830
rect 33310 7590 33400 7830
rect 33640 7590 33730 7830
rect 33970 7590 34060 7830
rect 34300 7590 34390 7830
rect 34630 7590 34720 7830
rect 34960 7590 35050 7830
rect 35290 7590 35430 7830
rect 28730 7500 35430 7590
rect 28730 7260 28780 7500
rect 29020 7260 29110 7500
rect 29350 7260 29440 7500
rect 29680 7260 29770 7500
rect 30010 7260 30100 7500
rect 30340 7260 30430 7500
rect 30670 7260 30760 7500
rect 31000 7260 31090 7500
rect 31330 7260 31420 7500
rect 31660 7260 31750 7500
rect 31990 7260 32080 7500
rect 32320 7260 32410 7500
rect 32650 7260 32740 7500
rect 32980 7260 33070 7500
rect 33310 7260 33400 7500
rect 33640 7260 33730 7500
rect 33970 7260 34060 7500
rect 34300 7260 34390 7500
rect 34630 7260 34720 7500
rect 34960 7260 35050 7500
rect 35290 7260 35430 7500
rect 28730 7170 35430 7260
rect 28730 6930 28780 7170
rect 29020 6930 29110 7170
rect 29350 6930 29440 7170
rect 29680 6930 29770 7170
rect 30010 6930 30100 7170
rect 30340 6930 30430 7170
rect 30670 6930 30760 7170
rect 31000 6930 31090 7170
rect 31330 6930 31420 7170
rect 31660 6930 31750 7170
rect 31990 6930 32080 7170
rect 32320 6930 32410 7170
rect 32650 6930 32740 7170
rect 32980 6930 33070 7170
rect 33310 6930 33400 7170
rect 33640 6930 33730 7170
rect 33970 6930 34060 7170
rect 34300 6930 34390 7170
rect 34630 6930 34720 7170
rect 34960 6930 35050 7170
rect 35290 6930 35430 7170
rect 28730 6840 35430 6930
rect 28730 6600 28780 6840
rect 29020 6600 29110 6840
rect 29350 6600 29440 6840
rect 29680 6600 29770 6840
rect 30010 6600 30100 6840
rect 30340 6600 30430 6840
rect 30670 6600 30760 6840
rect 31000 6600 31090 6840
rect 31330 6600 31420 6840
rect 31660 6600 31750 6840
rect 31990 6600 32080 6840
rect 32320 6600 32410 6840
rect 32650 6600 32740 6840
rect 32980 6600 33070 6840
rect 33310 6600 33400 6840
rect 33640 6600 33730 6840
rect 33970 6600 34060 6840
rect 34300 6600 34390 6840
rect 34630 6600 34720 6840
rect 34960 6600 35050 6840
rect 35290 6600 35430 6840
rect 28730 6510 35430 6600
rect 28730 6270 28780 6510
rect 29020 6270 29110 6510
rect 29350 6270 29440 6510
rect 29680 6270 29770 6510
rect 30010 6270 30100 6510
rect 30340 6270 30430 6510
rect 30670 6270 30760 6510
rect 31000 6270 31090 6510
rect 31330 6270 31420 6510
rect 31660 6270 31750 6510
rect 31990 6270 32080 6510
rect 32320 6270 32410 6510
rect 32650 6270 32740 6510
rect 32980 6270 33070 6510
rect 33310 6270 33400 6510
rect 33640 6270 33730 6510
rect 33970 6270 34060 6510
rect 34300 6270 34390 6510
rect 34630 6270 34720 6510
rect 34960 6270 35050 6510
rect 35290 6270 35430 6510
rect 28730 6180 35430 6270
rect 28730 5940 28780 6180
rect 29020 5940 29110 6180
rect 29350 5940 29440 6180
rect 29680 5940 29770 6180
rect 30010 5940 30100 6180
rect 30340 5940 30430 6180
rect 30670 5940 30760 6180
rect 31000 5940 31090 6180
rect 31330 5940 31420 6180
rect 31660 5940 31750 6180
rect 31990 5940 32080 6180
rect 32320 5940 32410 6180
rect 32650 5940 32740 6180
rect 32980 5940 33070 6180
rect 33310 5940 33400 6180
rect 33640 5940 33730 6180
rect 33970 5940 34060 6180
rect 34300 5940 34390 6180
rect 34630 5940 34720 6180
rect 34960 5940 35050 6180
rect 35290 5940 35430 6180
rect 28730 5850 35430 5940
rect 28730 5610 28780 5850
rect 29020 5610 29110 5850
rect 29350 5610 29440 5850
rect 29680 5610 29770 5850
rect 30010 5610 30100 5850
rect 30340 5610 30430 5850
rect 30670 5610 30760 5850
rect 31000 5610 31090 5850
rect 31330 5610 31420 5850
rect 31660 5610 31750 5850
rect 31990 5610 32080 5850
rect 32320 5610 32410 5850
rect 32650 5610 32740 5850
rect 32980 5610 33070 5850
rect 33310 5610 33400 5850
rect 33640 5610 33730 5850
rect 33970 5610 34060 5850
rect 34300 5610 34390 5850
rect 34630 5610 34720 5850
rect 34960 5610 35050 5850
rect 35290 5610 35430 5850
rect 28730 5520 35430 5610
rect 28730 5280 28780 5520
rect 29020 5280 29110 5520
rect 29350 5280 29440 5520
rect 29680 5280 29770 5520
rect 30010 5280 30100 5520
rect 30340 5280 30430 5520
rect 30670 5280 30760 5520
rect 31000 5280 31090 5520
rect 31330 5280 31420 5520
rect 31660 5280 31750 5520
rect 31990 5280 32080 5520
rect 32320 5280 32410 5520
rect 32650 5280 32740 5520
rect 32980 5280 33070 5520
rect 33310 5280 33400 5520
rect 33640 5280 33730 5520
rect 33970 5280 34060 5520
rect 34300 5280 34390 5520
rect 34630 5280 34720 5520
rect 34960 5280 35050 5520
rect 35290 5280 35430 5520
rect 28730 5190 35430 5280
rect 28730 4950 28780 5190
rect 29020 4950 29110 5190
rect 29350 4950 29440 5190
rect 29680 4950 29770 5190
rect 30010 4950 30100 5190
rect 30340 4950 30430 5190
rect 30670 4950 30760 5190
rect 31000 4950 31090 5190
rect 31330 4950 31420 5190
rect 31660 4950 31750 5190
rect 31990 4950 32080 5190
rect 32320 4950 32410 5190
rect 32650 4950 32740 5190
rect 32980 4950 33070 5190
rect 33310 4950 33400 5190
rect 33640 4950 33730 5190
rect 33970 4950 34060 5190
rect 34300 4950 34390 5190
rect 34630 4950 34720 5190
rect 34960 4950 35050 5190
rect 35290 4950 35430 5190
rect 28730 4860 35430 4950
rect 28730 4620 28780 4860
rect 29020 4620 29110 4860
rect 29350 4620 29440 4860
rect 29680 4620 29770 4860
rect 30010 4620 30100 4860
rect 30340 4620 30430 4860
rect 30670 4620 30760 4860
rect 31000 4620 31090 4860
rect 31330 4620 31420 4860
rect 31660 4620 31750 4860
rect 31990 4620 32080 4860
rect 32320 4620 32410 4860
rect 32650 4620 32740 4860
rect 32980 4620 33070 4860
rect 33310 4620 33400 4860
rect 33640 4620 33730 4860
rect 33970 4620 34060 4860
rect 34300 4620 34390 4860
rect 34630 4620 34720 4860
rect 34960 4620 35050 4860
rect 35290 4620 35430 4860
rect 28730 4530 35430 4620
rect 28730 4290 28780 4530
rect 29020 4290 29110 4530
rect 29350 4290 29440 4530
rect 29680 4290 29770 4530
rect 30010 4290 30100 4530
rect 30340 4290 30430 4530
rect 30670 4290 30760 4530
rect 31000 4290 31090 4530
rect 31330 4290 31420 4530
rect 31660 4290 31750 4530
rect 31990 4290 32080 4530
rect 32320 4290 32410 4530
rect 32650 4290 32740 4530
rect 32980 4290 33070 4530
rect 33310 4290 33400 4530
rect 33640 4290 33730 4530
rect 33970 4290 34060 4530
rect 34300 4290 34390 4530
rect 34630 4290 34720 4530
rect 34960 4290 35050 4530
rect 35290 4290 35430 4530
rect 28730 4200 35430 4290
rect 28730 3960 28780 4200
rect 29020 3960 29110 4200
rect 29350 3960 29440 4200
rect 29680 3960 29770 4200
rect 30010 3960 30100 4200
rect 30340 3960 30430 4200
rect 30670 3960 30760 4200
rect 31000 3960 31090 4200
rect 31330 3960 31420 4200
rect 31660 3960 31750 4200
rect 31990 3960 32080 4200
rect 32320 3960 32410 4200
rect 32650 3960 32740 4200
rect 32980 3960 33070 4200
rect 33310 3960 33400 4200
rect 33640 3960 33730 4200
rect 33970 3960 34060 4200
rect 34300 3960 34390 4200
rect 34630 3960 34720 4200
rect 34960 3960 35050 4200
rect 35290 3960 35430 4200
rect 28730 3870 35430 3960
rect 28730 3630 28780 3870
rect 29020 3630 29110 3870
rect 29350 3630 29440 3870
rect 29680 3630 29770 3870
rect 30010 3630 30100 3870
rect 30340 3630 30430 3870
rect 30670 3630 30760 3870
rect 31000 3630 31090 3870
rect 31330 3630 31420 3870
rect 31660 3630 31750 3870
rect 31990 3630 32080 3870
rect 32320 3630 32410 3870
rect 32650 3630 32740 3870
rect 32980 3630 33070 3870
rect 33310 3630 33400 3870
rect 33640 3630 33730 3870
rect 33970 3630 34060 3870
rect 34300 3630 34390 3870
rect 34630 3630 34720 3870
rect 34960 3630 35050 3870
rect 35290 3630 35430 3870
rect 28730 3540 35430 3630
rect 28730 3300 28780 3540
rect 29020 3300 29110 3540
rect 29350 3300 29440 3540
rect 29680 3300 29770 3540
rect 30010 3300 30100 3540
rect 30340 3300 30430 3540
rect 30670 3300 30760 3540
rect 31000 3300 31090 3540
rect 31330 3300 31420 3540
rect 31660 3300 31750 3540
rect 31990 3300 32080 3540
rect 32320 3300 32410 3540
rect 32650 3300 32740 3540
rect 32980 3300 33070 3540
rect 33310 3300 33400 3540
rect 33640 3300 33730 3540
rect 33970 3300 34060 3540
rect 34300 3300 34390 3540
rect 34630 3300 34720 3540
rect 34960 3300 35050 3540
rect 35290 3300 35430 3540
rect 28730 3210 35430 3300
rect 28730 2970 28780 3210
rect 29020 2970 29110 3210
rect 29350 2970 29440 3210
rect 29680 2970 29770 3210
rect 30010 2970 30100 3210
rect 30340 2970 30430 3210
rect 30670 2970 30760 3210
rect 31000 2970 31090 3210
rect 31330 2970 31420 3210
rect 31660 2970 31750 3210
rect 31990 2970 32080 3210
rect 32320 2970 32410 3210
rect 32650 2970 32740 3210
rect 32980 2970 33070 3210
rect 33310 2970 33400 3210
rect 33640 2970 33730 3210
rect 33970 2970 34060 3210
rect 34300 2970 34390 3210
rect 34630 2970 34720 3210
rect 34960 2970 35050 3210
rect 35290 2970 35430 3210
rect 28730 2880 35430 2970
rect 28730 2640 28780 2880
rect 29020 2640 29110 2880
rect 29350 2640 29440 2880
rect 29680 2640 29770 2880
rect 30010 2640 30100 2880
rect 30340 2640 30430 2880
rect 30670 2640 30760 2880
rect 31000 2640 31090 2880
rect 31330 2640 31420 2880
rect 31660 2640 31750 2880
rect 31990 2640 32080 2880
rect 32320 2640 32410 2880
rect 32650 2640 32740 2880
rect 32980 2640 33070 2880
rect 33310 2640 33400 2880
rect 33640 2640 33730 2880
rect 33970 2640 34060 2880
rect 34300 2640 34390 2880
rect 34630 2640 34720 2880
rect 34960 2640 35050 2880
rect 35290 2640 35430 2880
rect 28730 2550 35430 2640
rect 28730 2310 28780 2550
rect 29020 2310 29110 2550
rect 29350 2310 29440 2550
rect 29680 2310 29770 2550
rect 30010 2310 30100 2550
rect 30340 2310 30430 2550
rect 30670 2310 30760 2550
rect 31000 2310 31090 2550
rect 31330 2310 31420 2550
rect 31660 2310 31750 2550
rect 31990 2310 32080 2550
rect 32320 2310 32410 2550
rect 32650 2310 32740 2550
rect 32980 2310 33070 2550
rect 33310 2310 33400 2550
rect 33640 2310 33730 2550
rect 33970 2310 34060 2550
rect 34300 2310 34390 2550
rect 34630 2310 34720 2550
rect 34960 2310 35050 2550
rect 35290 2310 35430 2550
rect 28730 2220 35430 2310
rect 28730 1980 28780 2220
rect 29020 1980 29110 2220
rect 29350 1980 29440 2220
rect 29680 1980 29770 2220
rect 30010 1980 30100 2220
rect 30340 1980 30430 2220
rect 30670 1980 30760 2220
rect 31000 1980 31090 2220
rect 31330 1980 31420 2220
rect 31660 1980 31750 2220
rect 31990 1980 32080 2220
rect 32320 1980 32410 2220
rect 32650 1980 32740 2220
rect 32980 1980 33070 2220
rect 33310 1980 33400 2220
rect 33640 1980 33730 2220
rect 33970 1980 34060 2220
rect 34300 1980 34390 2220
rect 34630 1980 34720 2220
rect 34960 1980 35050 2220
rect 35290 1980 35430 2220
rect 28730 1890 35430 1980
rect 28730 1650 28780 1890
rect 29020 1650 29110 1890
rect 29350 1650 29440 1890
rect 29680 1650 29770 1890
rect 30010 1650 30100 1890
rect 30340 1650 30430 1890
rect 30670 1650 30760 1890
rect 31000 1650 31090 1890
rect 31330 1650 31420 1890
rect 31660 1650 31750 1890
rect 31990 1650 32080 1890
rect 32320 1650 32410 1890
rect 32650 1650 32740 1890
rect 32980 1650 33070 1890
rect 33310 1650 33400 1890
rect 33640 1650 33730 1890
rect 33970 1650 34060 1890
rect 34300 1650 34390 1890
rect 34630 1650 34720 1890
rect 34960 1650 35050 1890
rect 35290 1650 35430 1890
rect 28730 1560 35430 1650
rect 28730 1320 28780 1560
rect 29020 1320 29110 1560
rect 29350 1320 29440 1560
rect 29680 1320 29770 1560
rect 30010 1320 30100 1560
rect 30340 1320 30430 1560
rect 30670 1320 30760 1560
rect 31000 1320 31090 1560
rect 31330 1320 31420 1560
rect 31660 1320 31750 1560
rect 31990 1320 32080 1560
rect 32320 1320 32410 1560
rect 32650 1320 32740 1560
rect 32980 1320 33070 1560
rect 33310 1320 33400 1560
rect 33640 1320 33730 1560
rect 33970 1320 34060 1560
rect 34300 1320 34390 1560
rect 34630 1320 34720 1560
rect 34960 1320 35050 1560
rect 35290 1320 35430 1560
rect 28730 1180 35430 1320
rect 28730 230 35430 280
rect 28730 -10 28780 230
rect 29020 -10 29110 230
rect 29350 -10 29440 230
rect 29680 -10 29770 230
rect 30010 -10 30100 230
rect 30340 -10 30430 230
rect 30670 -10 30760 230
rect 31000 -10 31090 230
rect 31330 -10 31420 230
rect 31660 -10 31750 230
rect 31990 -10 32080 230
rect 32320 -10 32410 230
rect 32650 -10 32740 230
rect 32980 -10 33070 230
rect 33310 -10 33400 230
rect 33640 -10 33730 230
rect 33970 -10 34060 230
rect 34300 -10 34390 230
rect 34630 -10 34720 230
rect 34960 -10 35050 230
rect 35290 -10 35430 230
rect 28730 -100 35430 -10
rect 28730 -340 28780 -100
rect 29020 -340 29110 -100
rect 29350 -340 29440 -100
rect 29680 -340 29770 -100
rect 30010 -340 30100 -100
rect 30340 -340 30430 -100
rect 30670 -340 30760 -100
rect 31000 -340 31090 -100
rect 31330 -340 31420 -100
rect 31660 -340 31750 -100
rect 31990 -340 32080 -100
rect 32320 -340 32410 -100
rect 32650 -340 32740 -100
rect 32980 -340 33070 -100
rect 33310 -340 33400 -100
rect 33640 -340 33730 -100
rect 33970 -340 34060 -100
rect 34300 -340 34390 -100
rect 34630 -340 34720 -100
rect 34960 -340 35050 -100
rect 35290 -340 35430 -100
rect 28730 -430 35430 -340
rect 28730 -670 28780 -430
rect 29020 -670 29110 -430
rect 29350 -670 29440 -430
rect 29680 -670 29770 -430
rect 30010 -670 30100 -430
rect 30340 -670 30430 -430
rect 30670 -670 30760 -430
rect 31000 -670 31090 -430
rect 31330 -670 31420 -430
rect 31660 -670 31750 -430
rect 31990 -670 32080 -430
rect 32320 -670 32410 -430
rect 32650 -670 32740 -430
rect 32980 -670 33070 -430
rect 33310 -670 33400 -430
rect 33640 -670 33730 -430
rect 33970 -670 34060 -430
rect 34300 -670 34390 -430
rect 34630 -670 34720 -430
rect 34960 -670 35050 -430
rect 35290 -670 35430 -430
rect 28730 -760 35430 -670
rect 28730 -1000 28780 -760
rect 29020 -1000 29110 -760
rect 29350 -1000 29440 -760
rect 29680 -1000 29770 -760
rect 30010 -1000 30100 -760
rect 30340 -1000 30430 -760
rect 30670 -1000 30760 -760
rect 31000 -1000 31090 -760
rect 31330 -1000 31420 -760
rect 31660 -1000 31750 -760
rect 31990 -1000 32080 -760
rect 32320 -1000 32410 -760
rect 32650 -1000 32740 -760
rect 32980 -1000 33070 -760
rect 33310 -1000 33400 -760
rect 33640 -1000 33730 -760
rect 33970 -1000 34060 -760
rect 34300 -1000 34390 -760
rect 34630 -1000 34720 -760
rect 34960 -1000 35050 -760
rect 35290 -1000 35430 -760
rect 28730 -1090 35430 -1000
rect 28730 -1330 28780 -1090
rect 29020 -1330 29110 -1090
rect 29350 -1330 29440 -1090
rect 29680 -1330 29770 -1090
rect 30010 -1330 30100 -1090
rect 30340 -1330 30430 -1090
rect 30670 -1330 30760 -1090
rect 31000 -1330 31090 -1090
rect 31330 -1330 31420 -1090
rect 31660 -1330 31750 -1090
rect 31990 -1330 32080 -1090
rect 32320 -1330 32410 -1090
rect 32650 -1330 32740 -1090
rect 32980 -1330 33070 -1090
rect 33310 -1330 33400 -1090
rect 33640 -1330 33730 -1090
rect 33970 -1330 34060 -1090
rect 34300 -1330 34390 -1090
rect 34630 -1330 34720 -1090
rect 34960 -1330 35050 -1090
rect 35290 -1330 35430 -1090
rect 28730 -1420 35430 -1330
rect 28730 -1660 28780 -1420
rect 29020 -1660 29110 -1420
rect 29350 -1660 29440 -1420
rect 29680 -1660 29770 -1420
rect 30010 -1660 30100 -1420
rect 30340 -1660 30430 -1420
rect 30670 -1660 30760 -1420
rect 31000 -1660 31090 -1420
rect 31330 -1660 31420 -1420
rect 31660 -1660 31750 -1420
rect 31990 -1660 32080 -1420
rect 32320 -1660 32410 -1420
rect 32650 -1660 32740 -1420
rect 32980 -1660 33070 -1420
rect 33310 -1660 33400 -1420
rect 33640 -1660 33730 -1420
rect 33970 -1660 34060 -1420
rect 34300 -1660 34390 -1420
rect 34630 -1660 34720 -1420
rect 34960 -1660 35050 -1420
rect 35290 -1660 35430 -1420
rect 28730 -1750 35430 -1660
rect 28730 -1990 28780 -1750
rect 29020 -1990 29110 -1750
rect 29350 -1990 29440 -1750
rect 29680 -1990 29770 -1750
rect 30010 -1990 30100 -1750
rect 30340 -1990 30430 -1750
rect 30670 -1990 30760 -1750
rect 31000 -1990 31090 -1750
rect 31330 -1990 31420 -1750
rect 31660 -1990 31750 -1750
rect 31990 -1990 32080 -1750
rect 32320 -1990 32410 -1750
rect 32650 -1990 32740 -1750
rect 32980 -1990 33070 -1750
rect 33310 -1990 33400 -1750
rect 33640 -1990 33730 -1750
rect 33970 -1990 34060 -1750
rect 34300 -1990 34390 -1750
rect 34630 -1990 34720 -1750
rect 34960 -1990 35050 -1750
rect 35290 -1990 35430 -1750
rect 28730 -2080 35430 -1990
rect 28730 -2320 28780 -2080
rect 29020 -2320 29110 -2080
rect 29350 -2320 29440 -2080
rect 29680 -2320 29770 -2080
rect 30010 -2320 30100 -2080
rect 30340 -2320 30430 -2080
rect 30670 -2320 30760 -2080
rect 31000 -2320 31090 -2080
rect 31330 -2320 31420 -2080
rect 31660 -2320 31750 -2080
rect 31990 -2320 32080 -2080
rect 32320 -2320 32410 -2080
rect 32650 -2320 32740 -2080
rect 32980 -2320 33070 -2080
rect 33310 -2320 33400 -2080
rect 33640 -2320 33730 -2080
rect 33970 -2320 34060 -2080
rect 34300 -2320 34390 -2080
rect 34630 -2320 34720 -2080
rect 34960 -2320 35050 -2080
rect 35290 -2320 35430 -2080
rect 28730 -2410 35430 -2320
rect 28730 -2650 28780 -2410
rect 29020 -2650 29110 -2410
rect 29350 -2650 29440 -2410
rect 29680 -2650 29770 -2410
rect 30010 -2650 30100 -2410
rect 30340 -2650 30430 -2410
rect 30670 -2650 30760 -2410
rect 31000 -2650 31090 -2410
rect 31330 -2650 31420 -2410
rect 31660 -2650 31750 -2410
rect 31990 -2650 32080 -2410
rect 32320 -2650 32410 -2410
rect 32650 -2650 32740 -2410
rect 32980 -2650 33070 -2410
rect 33310 -2650 33400 -2410
rect 33640 -2650 33730 -2410
rect 33970 -2650 34060 -2410
rect 34300 -2650 34390 -2410
rect 34630 -2650 34720 -2410
rect 34960 -2650 35050 -2410
rect 35290 -2650 35430 -2410
rect 28730 -2740 35430 -2650
rect 28730 -2980 28780 -2740
rect 29020 -2980 29110 -2740
rect 29350 -2980 29440 -2740
rect 29680 -2980 29770 -2740
rect 30010 -2980 30100 -2740
rect 30340 -2980 30430 -2740
rect 30670 -2980 30760 -2740
rect 31000 -2980 31090 -2740
rect 31330 -2980 31420 -2740
rect 31660 -2980 31750 -2740
rect 31990 -2980 32080 -2740
rect 32320 -2980 32410 -2740
rect 32650 -2980 32740 -2740
rect 32980 -2980 33070 -2740
rect 33310 -2980 33400 -2740
rect 33640 -2980 33730 -2740
rect 33970 -2980 34060 -2740
rect 34300 -2980 34390 -2740
rect 34630 -2980 34720 -2740
rect 34960 -2980 35050 -2740
rect 35290 -2980 35430 -2740
rect 28730 -3070 35430 -2980
rect 28730 -3310 28780 -3070
rect 29020 -3310 29110 -3070
rect 29350 -3310 29440 -3070
rect 29680 -3310 29770 -3070
rect 30010 -3310 30100 -3070
rect 30340 -3310 30430 -3070
rect 30670 -3310 30760 -3070
rect 31000 -3310 31090 -3070
rect 31330 -3310 31420 -3070
rect 31660 -3310 31750 -3070
rect 31990 -3310 32080 -3070
rect 32320 -3310 32410 -3070
rect 32650 -3310 32740 -3070
rect 32980 -3310 33070 -3070
rect 33310 -3310 33400 -3070
rect 33640 -3310 33730 -3070
rect 33970 -3310 34060 -3070
rect 34300 -3310 34390 -3070
rect 34630 -3310 34720 -3070
rect 34960 -3310 35050 -3070
rect 35290 -3310 35430 -3070
rect 28730 -3400 35430 -3310
rect 28730 -3640 28780 -3400
rect 29020 -3640 29110 -3400
rect 29350 -3640 29440 -3400
rect 29680 -3640 29770 -3400
rect 30010 -3640 30100 -3400
rect 30340 -3640 30430 -3400
rect 30670 -3640 30760 -3400
rect 31000 -3640 31090 -3400
rect 31330 -3640 31420 -3400
rect 31660 -3640 31750 -3400
rect 31990 -3640 32080 -3400
rect 32320 -3640 32410 -3400
rect 32650 -3640 32740 -3400
rect 32980 -3640 33070 -3400
rect 33310 -3640 33400 -3400
rect 33640 -3640 33730 -3400
rect 33970 -3640 34060 -3400
rect 34300 -3640 34390 -3400
rect 34630 -3640 34720 -3400
rect 34960 -3640 35050 -3400
rect 35290 -3640 35430 -3400
rect 28730 -3730 35430 -3640
rect 28730 -3970 28780 -3730
rect 29020 -3970 29110 -3730
rect 29350 -3970 29440 -3730
rect 29680 -3970 29770 -3730
rect 30010 -3970 30100 -3730
rect 30340 -3970 30430 -3730
rect 30670 -3970 30760 -3730
rect 31000 -3970 31090 -3730
rect 31330 -3970 31420 -3730
rect 31660 -3970 31750 -3730
rect 31990 -3970 32080 -3730
rect 32320 -3970 32410 -3730
rect 32650 -3970 32740 -3730
rect 32980 -3970 33070 -3730
rect 33310 -3970 33400 -3730
rect 33640 -3970 33730 -3730
rect 33970 -3970 34060 -3730
rect 34300 -3970 34390 -3730
rect 34630 -3970 34720 -3730
rect 34960 -3970 35050 -3730
rect 35290 -3970 35430 -3730
rect 28730 -4060 35430 -3970
rect -1830 -4260 -280 -4080
rect -1830 -4500 -1650 -4260
rect -1410 -4500 -1320 -4260
rect -1080 -4500 -990 -4260
rect -750 -4500 -660 -4260
rect -420 -4500 -280 -4260
rect -1830 -4590 -280 -4500
rect -1830 -4830 -1650 -4590
rect -1410 -4830 -1320 -4590
rect -1080 -4830 -990 -4590
rect -750 -4830 -660 -4590
rect -420 -4830 -280 -4590
rect -1830 -4920 -280 -4830
rect -1830 -5160 -1650 -4920
rect -1410 -5160 -1320 -4920
rect -1080 -5160 -990 -4920
rect -750 -5160 -660 -4920
rect -420 -5160 -280 -4920
rect -1830 -5250 -280 -5160
rect -1830 -5490 -1650 -5250
rect -1410 -5490 -1320 -5250
rect -1080 -5490 -990 -5250
rect -750 -5490 -660 -5250
rect -420 -5490 -280 -5250
rect -1830 -5630 -280 -5490
rect 28730 -4300 28780 -4060
rect 29020 -4300 29110 -4060
rect 29350 -4300 29440 -4060
rect 29680 -4300 29770 -4060
rect 30010 -4300 30100 -4060
rect 30340 -4300 30430 -4060
rect 30670 -4300 30760 -4060
rect 31000 -4300 31090 -4060
rect 31330 -4300 31420 -4060
rect 31660 -4300 31750 -4060
rect 31990 -4300 32080 -4060
rect 32320 -4300 32410 -4060
rect 32650 -4300 32740 -4060
rect 32980 -4300 33070 -4060
rect 33310 -4300 33400 -4060
rect 33640 -4300 33730 -4060
rect 33970 -4300 34060 -4060
rect 34300 -4300 34390 -4060
rect 34630 -4300 34720 -4060
rect 34960 -4300 35050 -4060
rect 35290 -4300 35430 -4060
rect 28730 -4390 35430 -4300
rect 28730 -4630 28780 -4390
rect 29020 -4630 29110 -4390
rect 29350 -4630 29440 -4390
rect 29680 -4630 29770 -4390
rect 30010 -4630 30100 -4390
rect 30340 -4630 30430 -4390
rect 30670 -4630 30760 -4390
rect 31000 -4630 31090 -4390
rect 31330 -4630 31420 -4390
rect 31660 -4630 31750 -4390
rect 31990 -4630 32080 -4390
rect 32320 -4630 32410 -4390
rect 32650 -4630 32740 -4390
rect 32980 -4630 33070 -4390
rect 33310 -4630 33400 -4390
rect 33640 -4630 33730 -4390
rect 33970 -4630 34060 -4390
rect 34300 -4630 34390 -4390
rect 34630 -4630 34720 -4390
rect 34960 -4630 35050 -4390
rect 35290 -4630 35430 -4390
rect 28730 -4720 35430 -4630
rect 28730 -4960 28780 -4720
rect 29020 -4960 29110 -4720
rect 29350 -4960 29440 -4720
rect 29680 -4960 29770 -4720
rect 30010 -4960 30100 -4720
rect 30340 -4960 30430 -4720
rect 30670 -4960 30760 -4720
rect 31000 -4960 31090 -4720
rect 31330 -4960 31420 -4720
rect 31660 -4960 31750 -4720
rect 31990 -4960 32080 -4720
rect 32320 -4960 32410 -4720
rect 32650 -4960 32740 -4720
rect 32980 -4960 33070 -4720
rect 33310 -4960 33400 -4720
rect 33640 -4960 33730 -4720
rect 33970 -4960 34060 -4720
rect 34300 -4960 34390 -4720
rect 34630 -4960 34720 -4720
rect 34960 -4960 35050 -4720
rect 35290 -4960 35430 -4720
rect 28730 -5050 35430 -4960
rect 28730 -5290 28780 -5050
rect 29020 -5290 29110 -5050
rect 29350 -5290 29440 -5050
rect 29680 -5290 29770 -5050
rect 30010 -5290 30100 -5050
rect 30340 -5290 30430 -5050
rect 30670 -5290 30760 -5050
rect 31000 -5290 31090 -5050
rect 31330 -5290 31420 -5050
rect 31660 -5290 31750 -5050
rect 31990 -5290 32080 -5050
rect 32320 -5290 32410 -5050
rect 32650 -5290 32740 -5050
rect 32980 -5290 33070 -5050
rect 33310 -5290 33400 -5050
rect 33640 -5290 33730 -5050
rect 33970 -5290 34060 -5050
rect 34300 -5290 34390 -5050
rect 34630 -5290 34720 -5050
rect 34960 -5290 35050 -5050
rect 35290 -5290 35430 -5050
rect 28730 -5380 35430 -5290
rect 28730 -5620 28780 -5380
rect 29020 -5620 29110 -5380
rect 29350 -5620 29440 -5380
rect 29680 -5620 29770 -5380
rect 30010 -5620 30100 -5380
rect 30340 -5620 30430 -5380
rect 30670 -5620 30760 -5380
rect 31000 -5620 31090 -5380
rect 31330 -5620 31420 -5380
rect 31660 -5620 31750 -5380
rect 31990 -5620 32080 -5380
rect 32320 -5620 32410 -5380
rect 32650 -5620 32740 -5380
rect 32980 -5620 33070 -5380
rect 33310 -5620 33400 -5380
rect 33640 -5620 33730 -5380
rect 33970 -5620 34060 -5380
rect 34300 -5620 34390 -5380
rect 34630 -5620 34720 -5380
rect 34960 -5620 35050 -5380
rect 35290 -5620 35430 -5380
rect 28730 -5710 35430 -5620
rect 28730 -5950 28780 -5710
rect 29020 -5950 29110 -5710
rect 29350 -5950 29440 -5710
rect 29680 -5950 29770 -5710
rect 30010 -5950 30100 -5710
rect 30340 -5950 30430 -5710
rect 30670 -5950 30760 -5710
rect 31000 -5950 31090 -5710
rect 31330 -5950 31420 -5710
rect 31660 -5950 31750 -5710
rect 31990 -5950 32080 -5710
rect 32320 -5950 32410 -5710
rect 32650 -5950 32740 -5710
rect 32980 -5950 33070 -5710
rect 33310 -5950 33400 -5710
rect 33640 -5950 33730 -5710
rect 33970 -5950 34060 -5710
rect 34300 -5950 34390 -5710
rect 34630 -5950 34720 -5710
rect 34960 -5950 35050 -5710
rect 35290 -5950 35430 -5710
rect 28730 -6040 35430 -5950
rect 28730 -6280 28780 -6040
rect 29020 -6280 29110 -6040
rect 29350 -6280 29440 -6040
rect 29680 -6280 29770 -6040
rect 30010 -6280 30100 -6040
rect 30340 -6280 30430 -6040
rect 30670 -6280 30760 -6040
rect 31000 -6280 31090 -6040
rect 31330 -6280 31420 -6040
rect 31660 -6280 31750 -6040
rect 31990 -6280 32080 -6040
rect 32320 -6280 32410 -6040
rect 32650 -6280 32740 -6040
rect 32980 -6280 33070 -6040
rect 33310 -6280 33400 -6040
rect 33640 -6280 33730 -6040
rect 33970 -6280 34060 -6040
rect 34300 -6280 34390 -6040
rect 34630 -6280 34720 -6040
rect 34960 -6280 35050 -6040
rect 35290 -6280 35430 -6040
rect 28730 -6420 35430 -6280
rect -1830 -7660 -280 -7480
rect -1830 -7900 -1650 -7660
rect -1410 -7900 -1320 -7660
rect -1080 -7900 -990 -7660
rect -750 -7900 -660 -7660
rect -420 -7900 -280 -7660
rect -1830 -7990 -280 -7900
rect -1830 -8230 -1650 -7990
rect -1410 -8230 -1320 -7990
rect -1080 -8230 -990 -7990
rect -750 -8230 -660 -7990
rect -420 -8230 -280 -7990
rect -1830 -8320 -280 -8230
rect -1830 -8560 -1650 -8320
rect -1410 -8560 -1320 -8320
rect -1080 -8560 -990 -8320
rect -750 -8560 -660 -8320
rect -420 -8560 -280 -8320
rect -1830 -8650 -280 -8560
rect -1830 -8890 -1650 -8650
rect -1410 -8890 -1320 -8650
rect -1080 -8890 -990 -8650
rect -750 -8890 -660 -8650
rect -420 -8890 -280 -8650
rect -1830 -9030 -280 -8890
<< mimcap2contact >>
rect -4670 20550 -4430 20790
rect -4340 20550 -4100 20790
rect -4010 20550 -3770 20790
rect -3680 20550 -3440 20790
rect -3350 20550 -3110 20790
rect -3020 20550 -2780 20790
rect -2690 20550 -2450 20790
rect -2360 20550 -2120 20790
rect -2030 20550 -1790 20790
rect -1700 20550 -1460 20790
rect -1370 20550 -1130 20790
rect -1040 20550 -800 20790
rect -710 20550 -470 20790
rect -380 20550 -140 20790
rect -50 20550 190 20790
rect 280 20550 520 20790
rect 610 20550 850 20790
rect 940 20550 1180 20790
rect 1270 20550 1510 20790
rect 1600 20550 1840 20790
rect 1930 20550 2170 20790
rect 2260 20550 2500 20790
rect 2590 20550 2830 20790
rect 2920 20550 3160 20790
rect 3250 20550 3490 20790
rect 3580 20550 3820 20790
rect 3910 20550 4150 20790
rect 4240 20550 4480 20790
rect 4570 20550 4810 20790
rect 4900 20550 5140 20790
rect 5230 20550 5470 20790
rect 5560 20550 5800 20790
rect 5890 20550 6130 20790
rect 6220 20550 6460 20790
rect 6550 20550 6790 20790
rect 6880 20550 7120 20790
rect -4670 20220 -4430 20460
rect -4340 20220 -4100 20460
rect -4010 20220 -3770 20460
rect -3680 20220 -3440 20460
rect -3350 20220 -3110 20460
rect -3020 20220 -2780 20460
rect -2690 20220 -2450 20460
rect -2360 20220 -2120 20460
rect -2030 20220 -1790 20460
rect -1700 20220 -1460 20460
rect -1370 20220 -1130 20460
rect -1040 20220 -800 20460
rect -710 20220 -470 20460
rect -380 20220 -140 20460
rect -50 20220 190 20460
rect 280 20220 520 20460
rect 610 20220 850 20460
rect 940 20220 1180 20460
rect 1270 20220 1510 20460
rect 1600 20220 1840 20460
rect 1930 20220 2170 20460
rect 2260 20220 2500 20460
rect 2590 20220 2830 20460
rect 2920 20220 3160 20460
rect 3250 20220 3490 20460
rect 3580 20220 3820 20460
rect 3910 20220 4150 20460
rect 4240 20220 4480 20460
rect 4570 20220 4810 20460
rect 4900 20220 5140 20460
rect 5230 20220 5470 20460
rect 5560 20220 5800 20460
rect 5890 20220 6130 20460
rect 6220 20220 6460 20460
rect 6550 20220 6790 20460
rect 6880 20220 7120 20460
rect -4670 19890 -4430 20130
rect -4340 19890 -4100 20130
rect -4010 19890 -3770 20130
rect -3680 19890 -3440 20130
rect -3350 19890 -3110 20130
rect -3020 19890 -2780 20130
rect -2690 19890 -2450 20130
rect -2360 19890 -2120 20130
rect -2030 19890 -1790 20130
rect -1700 19890 -1460 20130
rect -1370 19890 -1130 20130
rect -1040 19890 -800 20130
rect -710 19890 -470 20130
rect -380 19890 -140 20130
rect -50 19890 190 20130
rect 280 19890 520 20130
rect 610 19890 850 20130
rect 940 19890 1180 20130
rect 1270 19890 1510 20130
rect 1600 19890 1840 20130
rect 1930 19890 2170 20130
rect 2260 19890 2500 20130
rect 2590 19890 2830 20130
rect 2920 19890 3160 20130
rect 3250 19890 3490 20130
rect 3580 19890 3820 20130
rect 3910 19890 4150 20130
rect 4240 19890 4480 20130
rect 4570 19890 4810 20130
rect 4900 19890 5140 20130
rect 5230 19890 5470 20130
rect 5560 19890 5800 20130
rect 5890 19890 6130 20130
rect 6220 19890 6460 20130
rect 6550 19890 6790 20130
rect 6880 19890 7120 20130
rect -4670 19560 -4430 19800
rect -4340 19560 -4100 19800
rect -4010 19560 -3770 19800
rect -3680 19560 -3440 19800
rect -3350 19560 -3110 19800
rect -3020 19560 -2780 19800
rect -2690 19560 -2450 19800
rect -2360 19560 -2120 19800
rect -2030 19560 -1790 19800
rect -1700 19560 -1460 19800
rect -1370 19560 -1130 19800
rect -1040 19560 -800 19800
rect -710 19560 -470 19800
rect -380 19560 -140 19800
rect -50 19560 190 19800
rect 280 19560 520 19800
rect 610 19560 850 19800
rect 940 19560 1180 19800
rect 1270 19560 1510 19800
rect 1600 19560 1840 19800
rect 1930 19560 2170 19800
rect 2260 19560 2500 19800
rect 2590 19560 2830 19800
rect 2920 19560 3160 19800
rect 3250 19560 3490 19800
rect 3580 19560 3820 19800
rect 3910 19560 4150 19800
rect 4240 19560 4480 19800
rect 4570 19560 4810 19800
rect 4900 19560 5140 19800
rect 5230 19560 5470 19800
rect 5560 19560 5800 19800
rect 5890 19560 6130 19800
rect 6220 19560 6460 19800
rect 6550 19560 6790 19800
rect 6880 19560 7120 19800
rect -4670 19230 -4430 19470
rect -4340 19230 -4100 19470
rect -4010 19230 -3770 19470
rect -3680 19230 -3440 19470
rect -3350 19230 -3110 19470
rect -3020 19230 -2780 19470
rect -2690 19230 -2450 19470
rect -2360 19230 -2120 19470
rect -2030 19230 -1790 19470
rect -1700 19230 -1460 19470
rect -1370 19230 -1130 19470
rect -1040 19230 -800 19470
rect -710 19230 -470 19470
rect -380 19230 -140 19470
rect -50 19230 190 19470
rect 280 19230 520 19470
rect 610 19230 850 19470
rect 940 19230 1180 19470
rect 1270 19230 1510 19470
rect 1600 19230 1840 19470
rect 1930 19230 2170 19470
rect 2260 19230 2500 19470
rect 2590 19230 2830 19470
rect 2920 19230 3160 19470
rect 3250 19230 3490 19470
rect 3580 19230 3820 19470
rect 3910 19230 4150 19470
rect 4240 19230 4480 19470
rect 4570 19230 4810 19470
rect 4900 19230 5140 19470
rect 5230 19230 5470 19470
rect 5560 19230 5800 19470
rect 5890 19230 6130 19470
rect 6220 19230 6460 19470
rect 6550 19230 6790 19470
rect 6880 19230 7120 19470
rect -4670 18900 -4430 19140
rect -4340 18900 -4100 19140
rect -4010 18900 -3770 19140
rect -3680 18900 -3440 19140
rect -3350 18900 -3110 19140
rect -3020 18900 -2780 19140
rect -2690 18900 -2450 19140
rect -2360 18900 -2120 19140
rect -2030 18900 -1790 19140
rect -1700 18900 -1460 19140
rect -1370 18900 -1130 19140
rect -1040 18900 -800 19140
rect -710 18900 -470 19140
rect -380 18900 -140 19140
rect -50 18900 190 19140
rect 280 18900 520 19140
rect 610 18900 850 19140
rect 940 18900 1180 19140
rect 1270 18900 1510 19140
rect 1600 18900 1840 19140
rect 1930 18900 2170 19140
rect 2260 18900 2500 19140
rect 2590 18900 2830 19140
rect 2920 18900 3160 19140
rect 3250 18900 3490 19140
rect 3580 18900 3820 19140
rect 3910 18900 4150 19140
rect 4240 18900 4480 19140
rect 4570 18900 4810 19140
rect 4900 18900 5140 19140
rect 5230 18900 5470 19140
rect 5560 18900 5800 19140
rect 5890 18900 6130 19140
rect 6220 18900 6460 19140
rect 6550 18900 6790 19140
rect 6880 18900 7120 19140
rect -4670 18570 -4430 18810
rect -4340 18570 -4100 18810
rect -4010 18570 -3770 18810
rect -3680 18570 -3440 18810
rect -3350 18570 -3110 18810
rect -3020 18570 -2780 18810
rect -2690 18570 -2450 18810
rect -2360 18570 -2120 18810
rect -2030 18570 -1790 18810
rect -1700 18570 -1460 18810
rect -1370 18570 -1130 18810
rect -1040 18570 -800 18810
rect -710 18570 -470 18810
rect -380 18570 -140 18810
rect -50 18570 190 18810
rect 280 18570 520 18810
rect 610 18570 850 18810
rect 940 18570 1180 18810
rect 1270 18570 1510 18810
rect 1600 18570 1840 18810
rect 1930 18570 2170 18810
rect 2260 18570 2500 18810
rect 2590 18570 2830 18810
rect 2920 18570 3160 18810
rect 3250 18570 3490 18810
rect 3580 18570 3820 18810
rect 3910 18570 4150 18810
rect 4240 18570 4480 18810
rect 4570 18570 4810 18810
rect 4900 18570 5140 18810
rect 5230 18570 5470 18810
rect 5560 18570 5800 18810
rect 5890 18570 6130 18810
rect 6220 18570 6460 18810
rect 6550 18570 6790 18810
rect 6880 18570 7120 18810
rect -4670 18240 -4430 18480
rect -4340 18240 -4100 18480
rect -4010 18240 -3770 18480
rect -3680 18240 -3440 18480
rect -3350 18240 -3110 18480
rect -3020 18240 -2780 18480
rect -2690 18240 -2450 18480
rect -2360 18240 -2120 18480
rect -2030 18240 -1790 18480
rect -1700 18240 -1460 18480
rect -1370 18240 -1130 18480
rect -1040 18240 -800 18480
rect -710 18240 -470 18480
rect -380 18240 -140 18480
rect -50 18240 190 18480
rect 280 18240 520 18480
rect 610 18240 850 18480
rect 940 18240 1180 18480
rect 1270 18240 1510 18480
rect 1600 18240 1840 18480
rect 1930 18240 2170 18480
rect 2260 18240 2500 18480
rect 2590 18240 2830 18480
rect 2920 18240 3160 18480
rect 3250 18240 3490 18480
rect 3580 18240 3820 18480
rect 3910 18240 4150 18480
rect 4240 18240 4480 18480
rect 4570 18240 4810 18480
rect 4900 18240 5140 18480
rect 5230 18240 5470 18480
rect 5560 18240 5800 18480
rect 5890 18240 6130 18480
rect 6220 18240 6460 18480
rect 6550 18240 6790 18480
rect 6880 18240 7120 18480
rect -4670 17910 -4430 18150
rect -4340 17910 -4100 18150
rect -4010 17910 -3770 18150
rect -3680 17910 -3440 18150
rect -3350 17910 -3110 18150
rect -3020 17910 -2780 18150
rect -2690 17910 -2450 18150
rect -2360 17910 -2120 18150
rect -2030 17910 -1790 18150
rect -1700 17910 -1460 18150
rect -1370 17910 -1130 18150
rect -1040 17910 -800 18150
rect -710 17910 -470 18150
rect -380 17910 -140 18150
rect -50 17910 190 18150
rect 280 17910 520 18150
rect 610 17910 850 18150
rect 940 17910 1180 18150
rect 1270 17910 1510 18150
rect 1600 17910 1840 18150
rect 1930 17910 2170 18150
rect 2260 17910 2500 18150
rect 2590 17910 2830 18150
rect 2920 17910 3160 18150
rect 3250 17910 3490 18150
rect 3580 17910 3820 18150
rect 3910 17910 4150 18150
rect 4240 17910 4480 18150
rect 4570 17910 4810 18150
rect 4900 17910 5140 18150
rect 5230 17910 5470 18150
rect 5560 17910 5800 18150
rect 5890 17910 6130 18150
rect 6220 17910 6460 18150
rect 6550 17910 6790 18150
rect 6880 17910 7120 18150
rect -4670 17580 -4430 17820
rect -4340 17580 -4100 17820
rect -4010 17580 -3770 17820
rect -3680 17580 -3440 17820
rect -3350 17580 -3110 17820
rect -3020 17580 -2780 17820
rect -2690 17580 -2450 17820
rect -2360 17580 -2120 17820
rect -2030 17580 -1790 17820
rect -1700 17580 -1460 17820
rect -1370 17580 -1130 17820
rect -1040 17580 -800 17820
rect -710 17580 -470 17820
rect -380 17580 -140 17820
rect -50 17580 190 17820
rect 280 17580 520 17820
rect 610 17580 850 17820
rect 940 17580 1180 17820
rect 1270 17580 1510 17820
rect 1600 17580 1840 17820
rect 1930 17580 2170 17820
rect 2260 17580 2500 17820
rect 2590 17580 2830 17820
rect 2920 17580 3160 17820
rect 3250 17580 3490 17820
rect 3580 17580 3820 17820
rect 3910 17580 4150 17820
rect 4240 17580 4480 17820
rect 4570 17580 4810 17820
rect 4900 17580 5140 17820
rect 5230 17580 5470 17820
rect 5560 17580 5800 17820
rect 5890 17580 6130 17820
rect 6220 17580 6460 17820
rect 6550 17580 6790 17820
rect 6880 17580 7120 17820
rect -4670 17250 -4430 17490
rect -4340 17250 -4100 17490
rect -4010 17250 -3770 17490
rect -3680 17250 -3440 17490
rect -3350 17250 -3110 17490
rect -3020 17250 -2780 17490
rect -2690 17250 -2450 17490
rect -2360 17250 -2120 17490
rect -2030 17250 -1790 17490
rect -1700 17250 -1460 17490
rect -1370 17250 -1130 17490
rect -1040 17250 -800 17490
rect -710 17250 -470 17490
rect -380 17250 -140 17490
rect -50 17250 190 17490
rect 280 17250 520 17490
rect 610 17250 850 17490
rect 940 17250 1180 17490
rect 1270 17250 1510 17490
rect 1600 17250 1840 17490
rect 1930 17250 2170 17490
rect 2260 17250 2500 17490
rect 2590 17250 2830 17490
rect 2920 17250 3160 17490
rect 3250 17250 3490 17490
rect 3580 17250 3820 17490
rect 3910 17250 4150 17490
rect 4240 17250 4480 17490
rect 4570 17250 4810 17490
rect 4900 17250 5140 17490
rect 5230 17250 5470 17490
rect 5560 17250 5800 17490
rect 5890 17250 6130 17490
rect 6220 17250 6460 17490
rect 6550 17250 6790 17490
rect 6880 17250 7120 17490
rect -4670 16920 -4430 17160
rect -4340 16920 -4100 17160
rect -4010 16920 -3770 17160
rect -3680 16920 -3440 17160
rect -3350 16920 -3110 17160
rect -3020 16920 -2780 17160
rect -2690 16920 -2450 17160
rect -2360 16920 -2120 17160
rect -2030 16920 -1790 17160
rect -1700 16920 -1460 17160
rect -1370 16920 -1130 17160
rect -1040 16920 -800 17160
rect -710 16920 -470 17160
rect -380 16920 -140 17160
rect -50 16920 190 17160
rect 280 16920 520 17160
rect 610 16920 850 17160
rect 940 16920 1180 17160
rect 1270 16920 1510 17160
rect 1600 16920 1840 17160
rect 1930 16920 2170 17160
rect 2260 16920 2500 17160
rect 2590 16920 2830 17160
rect 2920 16920 3160 17160
rect 3250 16920 3490 17160
rect 3580 16920 3820 17160
rect 3910 16920 4150 17160
rect 4240 16920 4480 17160
rect 4570 16920 4810 17160
rect 4900 16920 5140 17160
rect 5230 16920 5470 17160
rect 5560 16920 5800 17160
rect 5890 16920 6130 17160
rect 6220 16920 6460 17160
rect 6550 16920 6790 17160
rect 6880 16920 7120 17160
rect -4670 16590 -4430 16830
rect -4340 16590 -4100 16830
rect -4010 16590 -3770 16830
rect -3680 16590 -3440 16830
rect -3350 16590 -3110 16830
rect -3020 16590 -2780 16830
rect -2690 16590 -2450 16830
rect -2360 16590 -2120 16830
rect -2030 16590 -1790 16830
rect -1700 16590 -1460 16830
rect -1370 16590 -1130 16830
rect -1040 16590 -800 16830
rect -710 16590 -470 16830
rect -380 16590 -140 16830
rect -50 16590 190 16830
rect 280 16590 520 16830
rect 610 16590 850 16830
rect 940 16590 1180 16830
rect 1270 16590 1510 16830
rect 1600 16590 1840 16830
rect 1930 16590 2170 16830
rect 2260 16590 2500 16830
rect 2590 16590 2830 16830
rect 2920 16590 3160 16830
rect 3250 16590 3490 16830
rect 3580 16590 3820 16830
rect 3910 16590 4150 16830
rect 4240 16590 4480 16830
rect 4570 16590 4810 16830
rect 4900 16590 5140 16830
rect 5230 16590 5470 16830
rect 5560 16590 5800 16830
rect 5890 16590 6130 16830
rect 6220 16590 6460 16830
rect 6550 16590 6790 16830
rect 6880 16590 7120 16830
rect -4670 16260 -4430 16500
rect -4340 16260 -4100 16500
rect -4010 16260 -3770 16500
rect -3680 16260 -3440 16500
rect -3350 16260 -3110 16500
rect -3020 16260 -2780 16500
rect -2690 16260 -2450 16500
rect -2360 16260 -2120 16500
rect -2030 16260 -1790 16500
rect -1700 16260 -1460 16500
rect -1370 16260 -1130 16500
rect -1040 16260 -800 16500
rect -710 16260 -470 16500
rect -380 16260 -140 16500
rect -50 16260 190 16500
rect 280 16260 520 16500
rect 610 16260 850 16500
rect 940 16260 1180 16500
rect 1270 16260 1510 16500
rect 1600 16260 1840 16500
rect 1930 16260 2170 16500
rect 2260 16260 2500 16500
rect 2590 16260 2830 16500
rect 2920 16260 3160 16500
rect 3250 16260 3490 16500
rect 3580 16260 3820 16500
rect 3910 16260 4150 16500
rect 4240 16260 4480 16500
rect 4570 16260 4810 16500
rect 4900 16260 5140 16500
rect 5230 16260 5470 16500
rect 5560 16260 5800 16500
rect 5890 16260 6130 16500
rect 6220 16260 6460 16500
rect 6550 16260 6790 16500
rect 6880 16260 7120 16500
rect -4670 15930 -4430 16170
rect -4340 15930 -4100 16170
rect -4010 15930 -3770 16170
rect -3680 15930 -3440 16170
rect -3350 15930 -3110 16170
rect -3020 15930 -2780 16170
rect -2690 15930 -2450 16170
rect -2360 15930 -2120 16170
rect -2030 15930 -1790 16170
rect -1700 15930 -1460 16170
rect -1370 15930 -1130 16170
rect -1040 15930 -800 16170
rect -710 15930 -470 16170
rect -380 15930 -140 16170
rect -50 15930 190 16170
rect 280 15930 520 16170
rect 610 15930 850 16170
rect 940 15930 1180 16170
rect 1270 15930 1510 16170
rect 1600 15930 1840 16170
rect 1930 15930 2170 16170
rect 2260 15930 2500 16170
rect 2590 15930 2830 16170
rect 2920 15930 3160 16170
rect 3250 15930 3490 16170
rect 3580 15930 3820 16170
rect 3910 15930 4150 16170
rect 4240 15930 4480 16170
rect 4570 15930 4810 16170
rect 4900 15930 5140 16170
rect 5230 15930 5470 16170
rect 5560 15930 5800 16170
rect 5890 15930 6130 16170
rect 6220 15930 6460 16170
rect 6550 15930 6790 16170
rect 6880 15930 7120 16170
rect -4670 15600 -4430 15840
rect -4340 15600 -4100 15840
rect -4010 15600 -3770 15840
rect -3680 15600 -3440 15840
rect -3350 15600 -3110 15840
rect -3020 15600 -2780 15840
rect -2690 15600 -2450 15840
rect -2360 15600 -2120 15840
rect -2030 15600 -1790 15840
rect -1700 15600 -1460 15840
rect -1370 15600 -1130 15840
rect -1040 15600 -800 15840
rect -710 15600 -470 15840
rect -380 15600 -140 15840
rect -50 15600 190 15840
rect 280 15600 520 15840
rect 610 15600 850 15840
rect 940 15600 1180 15840
rect 1270 15600 1510 15840
rect 1600 15600 1840 15840
rect 1930 15600 2170 15840
rect 2260 15600 2500 15840
rect 2590 15600 2830 15840
rect 2920 15600 3160 15840
rect 3250 15600 3490 15840
rect 3580 15600 3820 15840
rect 3910 15600 4150 15840
rect 4240 15600 4480 15840
rect 4570 15600 4810 15840
rect 4900 15600 5140 15840
rect 5230 15600 5470 15840
rect 5560 15600 5800 15840
rect 5890 15600 6130 15840
rect 6220 15600 6460 15840
rect 6550 15600 6790 15840
rect 6880 15600 7120 15840
rect -4670 15270 -4430 15510
rect -4340 15270 -4100 15510
rect -4010 15270 -3770 15510
rect -3680 15270 -3440 15510
rect -3350 15270 -3110 15510
rect -3020 15270 -2780 15510
rect -2690 15270 -2450 15510
rect -2360 15270 -2120 15510
rect -2030 15270 -1790 15510
rect -1700 15270 -1460 15510
rect -1370 15270 -1130 15510
rect -1040 15270 -800 15510
rect -710 15270 -470 15510
rect -380 15270 -140 15510
rect -50 15270 190 15510
rect 280 15270 520 15510
rect 610 15270 850 15510
rect 940 15270 1180 15510
rect 1270 15270 1510 15510
rect 1600 15270 1840 15510
rect 1930 15270 2170 15510
rect 2260 15270 2500 15510
rect 2590 15270 2830 15510
rect 2920 15270 3160 15510
rect 3250 15270 3490 15510
rect 3580 15270 3820 15510
rect 3910 15270 4150 15510
rect 4240 15270 4480 15510
rect 4570 15270 4810 15510
rect 4900 15270 5140 15510
rect 5230 15270 5470 15510
rect 5560 15270 5800 15510
rect 5890 15270 6130 15510
rect 6220 15270 6460 15510
rect 6550 15270 6790 15510
rect 6880 15270 7120 15510
rect -4670 14940 -4430 15180
rect -4340 14940 -4100 15180
rect -4010 14940 -3770 15180
rect -3680 14940 -3440 15180
rect -3350 14940 -3110 15180
rect -3020 14940 -2780 15180
rect -2690 14940 -2450 15180
rect -2360 14940 -2120 15180
rect -2030 14940 -1790 15180
rect -1700 14940 -1460 15180
rect -1370 14940 -1130 15180
rect -1040 14940 -800 15180
rect -710 14940 -470 15180
rect -380 14940 -140 15180
rect -50 14940 190 15180
rect 280 14940 520 15180
rect 610 14940 850 15180
rect 940 14940 1180 15180
rect 1270 14940 1510 15180
rect 1600 14940 1840 15180
rect 1930 14940 2170 15180
rect 2260 14940 2500 15180
rect 2590 14940 2830 15180
rect 2920 14940 3160 15180
rect 3250 14940 3490 15180
rect 3580 14940 3820 15180
rect 3910 14940 4150 15180
rect 4240 14940 4480 15180
rect 4570 14940 4810 15180
rect 4900 14940 5140 15180
rect 5230 14940 5470 15180
rect 5560 14940 5800 15180
rect 5890 14940 6130 15180
rect 6220 14940 6460 15180
rect 6550 14940 6790 15180
rect 6880 14940 7120 15180
rect -4670 14610 -4430 14850
rect -4340 14610 -4100 14850
rect -4010 14610 -3770 14850
rect -3680 14610 -3440 14850
rect -3350 14610 -3110 14850
rect -3020 14610 -2780 14850
rect -2690 14610 -2450 14850
rect -2360 14610 -2120 14850
rect -2030 14610 -1790 14850
rect -1700 14610 -1460 14850
rect -1370 14610 -1130 14850
rect -1040 14610 -800 14850
rect -710 14610 -470 14850
rect -380 14610 -140 14850
rect -50 14610 190 14850
rect 280 14610 520 14850
rect 610 14610 850 14850
rect 940 14610 1180 14850
rect 1270 14610 1510 14850
rect 1600 14610 1840 14850
rect 1930 14610 2170 14850
rect 2260 14610 2500 14850
rect 2590 14610 2830 14850
rect 2920 14610 3160 14850
rect 3250 14610 3490 14850
rect 3580 14610 3820 14850
rect 3910 14610 4150 14850
rect 4240 14610 4480 14850
rect 4570 14610 4810 14850
rect 4900 14610 5140 14850
rect 5230 14610 5470 14850
rect 5560 14610 5800 14850
rect 5890 14610 6130 14850
rect 6220 14610 6460 14850
rect 6550 14610 6790 14850
rect 6880 14610 7120 14850
rect -4670 14280 -4430 14520
rect -4340 14280 -4100 14520
rect -4010 14280 -3770 14520
rect -3680 14280 -3440 14520
rect -3350 14280 -3110 14520
rect -3020 14280 -2780 14520
rect -2690 14280 -2450 14520
rect -2360 14280 -2120 14520
rect -2030 14280 -1790 14520
rect -1700 14280 -1460 14520
rect -1370 14280 -1130 14520
rect -1040 14280 -800 14520
rect -710 14280 -470 14520
rect -380 14280 -140 14520
rect -50 14280 190 14520
rect 280 14280 520 14520
rect 610 14280 850 14520
rect 940 14280 1180 14520
rect 1270 14280 1510 14520
rect 1600 14280 1840 14520
rect 1930 14280 2170 14520
rect 2260 14280 2500 14520
rect 2590 14280 2830 14520
rect 2920 14280 3160 14520
rect 3250 14280 3490 14520
rect 3580 14280 3820 14520
rect 3910 14280 4150 14520
rect 4240 14280 4480 14520
rect 4570 14280 4810 14520
rect 4900 14280 5140 14520
rect 5230 14280 5470 14520
rect 5560 14280 5800 14520
rect 5890 14280 6130 14520
rect 6220 14280 6460 14520
rect 6550 14280 6790 14520
rect 6880 14280 7120 14520
rect -4670 13950 -4430 14190
rect -4340 13950 -4100 14190
rect -4010 13950 -3770 14190
rect -3680 13950 -3440 14190
rect -3350 13950 -3110 14190
rect -3020 13950 -2780 14190
rect -2690 13950 -2450 14190
rect -2360 13950 -2120 14190
rect -2030 13950 -1790 14190
rect -1700 13950 -1460 14190
rect -1370 13950 -1130 14190
rect -1040 13950 -800 14190
rect -710 13950 -470 14190
rect -380 13950 -140 14190
rect -50 13950 190 14190
rect 280 13950 520 14190
rect 610 13950 850 14190
rect 940 13950 1180 14190
rect 1270 13950 1510 14190
rect 1600 13950 1840 14190
rect 1930 13950 2170 14190
rect 2260 13950 2500 14190
rect 2590 13950 2830 14190
rect 2920 13950 3160 14190
rect 3250 13950 3490 14190
rect 3580 13950 3820 14190
rect 3910 13950 4150 14190
rect 4240 13950 4480 14190
rect 4570 13950 4810 14190
rect 4900 13950 5140 14190
rect 5230 13950 5470 14190
rect 5560 13950 5800 14190
rect 5890 13950 6130 14190
rect 6220 13950 6460 14190
rect 6550 13950 6790 14190
rect 6880 13950 7120 14190
rect -4670 13620 -4430 13860
rect -4340 13620 -4100 13860
rect -4010 13620 -3770 13860
rect -3680 13620 -3440 13860
rect -3350 13620 -3110 13860
rect -3020 13620 -2780 13860
rect -2690 13620 -2450 13860
rect -2360 13620 -2120 13860
rect -2030 13620 -1790 13860
rect -1700 13620 -1460 13860
rect -1370 13620 -1130 13860
rect -1040 13620 -800 13860
rect -710 13620 -470 13860
rect -380 13620 -140 13860
rect -50 13620 190 13860
rect 280 13620 520 13860
rect 610 13620 850 13860
rect 940 13620 1180 13860
rect 1270 13620 1510 13860
rect 1600 13620 1840 13860
rect 1930 13620 2170 13860
rect 2260 13620 2500 13860
rect 2590 13620 2830 13860
rect 2920 13620 3160 13860
rect 3250 13620 3490 13860
rect 3580 13620 3820 13860
rect 3910 13620 4150 13860
rect 4240 13620 4480 13860
rect 4570 13620 4810 13860
rect 4900 13620 5140 13860
rect 5230 13620 5470 13860
rect 5560 13620 5800 13860
rect 5890 13620 6130 13860
rect 6220 13620 6460 13860
rect 6550 13620 6790 13860
rect 6880 13620 7120 13860
rect -4670 13290 -4430 13530
rect -4340 13290 -4100 13530
rect -4010 13290 -3770 13530
rect -3680 13290 -3440 13530
rect -3350 13290 -3110 13530
rect -3020 13290 -2780 13530
rect -2690 13290 -2450 13530
rect -2360 13290 -2120 13530
rect -2030 13290 -1790 13530
rect -1700 13290 -1460 13530
rect -1370 13290 -1130 13530
rect -1040 13290 -800 13530
rect -710 13290 -470 13530
rect -380 13290 -140 13530
rect -50 13290 190 13530
rect 280 13290 520 13530
rect 610 13290 850 13530
rect 940 13290 1180 13530
rect 1270 13290 1510 13530
rect 1600 13290 1840 13530
rect 1930 13290 2170 13530
rect 2260 13290 2500 13530
rect 2590 13290 2830 13530
rect 2920 13290 3160 13530
rect 3250 13290 3490 13530
rect 3580 13290 3820 13530
rect 3910 13290 4150 13530
rect 4240 13290 4480 13530
rect 4570 13290 4810 13530
rect 4900 13290 5140 13530
rect 5230 13290 5470 13530
rect 5560 13290 5800 13530
rect 5890 13290 6130 13530
rect 6220 13290 6460 13530
rect 6550 13290 6790 13530
rect 6880 13290 7120 13530
rect -4670 12960 -4430 13200
rect -4340 12960 -4100 13200
rect -4010 12960 -3770 13200
rect -3680 12960 -3440 13200
rect -3350 12960 -3110 13200
rect -3020 12960 -2780 13200
rect -2690 12960 -2450 13200
rect -2360 12960 -2120 13200
rect -2030 12960 -1790 13200
rect -1700 12960 -1460 13200
rect -1370 12960 -1130 13200
rect -1040 12960 -800 13200
rect -710 12960 -470 13200
rect -380 12960 -140 13200
rect -50 12960 190 13200
rect 280 12960 520 13200
rect 610 12960 850 13200
rect 940 12960 1180 13200
rect 1270 12960 1510 13200
rect 1600 12960 1840 13200
rect 1930 12960 2170 13200
rect 2260 12960 2500 13200
rect 2590 12960 2830 13200
rect 2920 12960 3160 13200
rect 3250 12960 3490 13200
rect 3580 12960 3820 13200
rect 3910 12960 4150 13200
rect 4240 12960 4480 13200
rect 4570 12960 4810 13200
rect 4900 12960 5140 13200
rect 5230 12960 5470 13200
rect 5560 12960 5800 13200
rect 5890 12960 6130 13200
rect 6220 12960 6460 13200
rect 6550 12960 6790 13200
rect 6880 12960 7120 13200
rect -4670 12630 -4430 12870
rect -4340 12630 -4100 12870
rect -4010 12630 -3770 12870
rect -3680 12630 -3440 12870
rect -3350 12630 -3110 12870
rect -3020 12630 -2780 12870
rect -2690 12630 -2450 12870
rect -2360 12630 -2120 12870
rect -2030 12630 -1790 12870
rect -1700 12630 -1460 12870
rect -1370 12630 -1130 12870
rect -1040 12630 -800 12870
rect -710 12630 -470 12870
rect -380 12630 -140 12870
rect -50 12630 190 12870
rect 280 12630 520 12870
rect 610 12630 850 12870
rect 940 12630 1180 12870
rect 1270 12630 1510 12870
rect 1600 12630 1840 12870
rect 1930 12630 2170 12870
rect 2260 12630 2500 12870
rect 2590 12630 2830 12870
rect 2920 12630 3160 12870
rect 3250 12630 3490 12870
rect 3580 12630 3820 12870
rect 3910 12630 4150 12870
rect 4240 12630 4480 12870
rect 4570 12630 4810 12870
rect 4900 12630 5140 12870
rect 5230 12630 5470 12870
rect 5560 12630 5800 12870
rect 5890 12630 6130 12870
rect 6220 12630 6460 12870
rect 6550 12630 6790 12870
rect 6880 12630 7120 12870
rect -4670 12300 -4430 12540
rect -4340 12300 -4100 12540
rect -4010 12300 -3770 12540
rect -3680 12300 -3440 12540
rect -3350 12300 -3110 12540
rect -3020 12300 -2780 12540
rect -2690 12300 -2450 12540
rect -2360 12300 -2120 12540
rect -2030 12300 -1790 12540
rect -1700 12300 -1460 12540
rect -1370 12300 -1130 12540
rect -1040 12300 -800 12540
rect -710 12300 -470 12540
rect -380 12300 -140 12540
rect -50 12300 190 12540
rect 280 12300 520 12540
rect 610 12300 850 12540
rect 940 12300 1180 12540
rect 1270 12300 1510 12540
rect 1600 12300 1840 12540
rect 1930 12300 2170 12540
rect 2260 12300 2500 12540
rect 2590 12300 2830 12540
rect 2920 12300 3160 12540
rect 3250 12300 3490 12540
rect 3580 12300 3820 12540
rect 3910 12300 4150 12540
rect 4240 12300 4480 12540
rect 4570 12300 4810 12540
rect 4900 12300 5140 12540
rect 5230 12300 5470 12540
rect 5560 12300 5800 12540
rect 5890 12300 6130 12540
rect 6220 12300 6460 12540
rect 6550 12300 6790 12540
rect 6880 12300 7120 12540
rect -4670 11970 -4430 12210
rect -4340 11970 -4100 12210
rect -4010 11970 -3770 12210
rect -3680 11970 -3440 12210
rect -3350 11970 -3110 12210
rect -3020 11970 -2780 12210
rect -2690 11970 -2450 12210
rect -2360 11970 -2120 12210
rect -2030 11970 -1790 12210
rect -1700 11970 -1460 12210
rect -1370 11970 -1130 12210
rect -1040 11970 -800 12210
rect -710 11970 -470 12210
rect -380 11970 -140 12210
rect -50 11970 190 12210
rect 280 11970 520 12210
rect 610 11970 850 12210
rect 940 11970 1180 12210
rect 1270 11970 1510 12210
rect 1600 11970 1840 12210
rect 1930 11970 2170 12210
rect 2260 11970 2500 12210
rect 2590 11970 2830 12210
rect 2920 11970 3160 12210
rect 3250 11970 3490 12210
rect 3580 11970 3820 12210
rect 3910 11970 4150 12210
rect 4240 11970 4480 12210
rect 4570 11970 4810 12210
rect 4900 11970 5140 12210
rect 5230 11970 5470 12210
rect 5560 11970 5800 12210
rect 5890 11970 6130 12210
rect 6220 11970 6460 12210
rect 6550 11970 6790 12210
rect 6880 11970 7120 12210
rect -4670 11640 -4430 11880
rect -4340 11640 -4100 11880
rect -4010 11640 -3770 11880
rect -3680 11640 -3440 11880
rect -3350 11640 -3110 11880
rect -3020 11640 -2780 11880
rect -2690 11640 -2450 11880
rect -2360 11640 -2120 11880
rect -2030 11640 -1790 11880
rect -1700 11640 -1460 11880
rect -1370 11640 -1130 11880
rect -1040 11640 -800 11880
rect -710 11640 -470 11880
rect -380 11640 -140 11880
rect -50 11640 190 11880
rect 280 11640 520 11880
rect 610 11640 850 11880
rect 940 11640 1180 11880
rect 1270 11640 1510 11880
rect 1600 11640 1840 11880
rect 1930 11640 2170 11880
rect 2260 11640 2500 11880
rect 2590 11640 2830 11880
rect 2920 11640 3160 11880
rect 3250 11640 3490 11880
rect 3580 11640 3820 11880
rect 3910 11640 4150 11880
rect 4240 11640 4480 11880
rect 4570 11640 4810 11880
rect 4900 11640 5140 11880
rect 5230 11640 5470 11880
rect 5560 11640 5800 11880
rect 5890 11640 6130 11880
rect 6220 11640 6460 11880
rect 6550 11640 6790 11880
rect 6880 11640 7120 11880
rect -4670 11310 -4430 11550
rect -4340 11310 -4100 11550
rect -4010 11310 -3770 11550
rect -3680 11310 -3440 11550
rect -3350 11310 -3110 11550
rect -3020 11310 -2780 11550
rect -2690 11310 -2450 11550
rect -2360 11310 -2120 11550
rect -2030 11310 -1790 11550
rect -1700 11310 -1460 11550
rect -1370 11310 -1130 11550
rect -1040 11310 -800 11550
rect -710 11310 -470 11550
rect -380 11310 -140 11550
rect -50 11310 190 11550
rect 280 11310 520 11550
rect 610 11310 850 11550
rect 940 11310 1180 11550
rect 1270 11310 1510 11550
rect 1600 11310 1840 11550
rect 1930 11310 2170 11550
rect 2260 11310 2500 11550
rect 2590 11310 2830 11550
rect 2920 11310 3160 11550
rect 3250 11310 3490 11550
rect 3580 11310 3820 11550
rect 3910 11310 4150 11550
rect 4240 11310 4480 11550
rect 4570 11310 4810 11550
rect 4900 11310 5140 11550
rect 5230 11310 5470 11550
rect 5560 11310 5800 11550
rect 5890 11310 6130 11550
rect 6220 11310 6460 11550
rect 6550 11310 6790 11550
rect 6880 11310 7120 11550
rect -4670 10980 -4430 11220
rect -4340 10980 -4100 11220
rect -4010 10980 -3770 11220
rect -3680 10980 -3440 11220
rect -3350 10980 -3110 11220
rect -3020 10980 -2780 11220
rect -2690 10980 -2450 11220
rect -2360 10980 -2120 11220
rect -2030 10980 -1790 11220
rect -1700 10980 -1460 11220
rect -1370 10980 -1130 11220
rect -1040 10980 -800 11220
rect -710 10980 -470 11220
rect -380 10980 -140 11220
rect -50 10980 190 11220
rect 280 10980 520 11220
rect 610 10980 850 11220
rect 940 10980 1180 11220
rect 1270 10980 1510 11220
rect 1600 10980 1840 11220
rect 1930 10980 2170 11220
rect 2260 10980 2500 11220
rect 2590 10980 2830 11220
rect 2920 10980 3160 11220
rect 3250 10980 3490 11220
rect 3580 10980 3820 11220
rect 3910 10980 4150 11220
rect 4240 10980 4480 11220
rect 4570 10980 4810 11220
rect 4900 10980 5140 11220
rect 5230 10980 5470 11220
rect 5560 10980 5800 11220
rect 5890 10980 6130 11220
rect 6220 10980 6460 11220
rect 6550 10980 6790 11220
rect 6880 10980 7120 11220
rect -4670 10650 -4430 10890
rect -4340 10650 -4100 10890
rect -4010 10650 -3770 10890
rect -3680 10650 -3440 10890
rect -3350 10650 -3110 10890
rect -3020 10650 -2780 10890
rect -2690 10650 -2450 10890
rect -2360 10650 -2120 10890
rect -2030 10650 -1790 10890
rect -1700 10650 -1460 10890
rect -1370 10650 -1130 10890
rect -1040 10650 -800 10890
rect -710 10650 -470 10890
rect -380 10650 -140 10890
rect -50 10650 190 10890
rect 280 10650 520 10890
rect 610 10650 850 10890
rect 940 10650 1180 10890
rect 1270 10650 1510 10890
rect 1600 10650 1840 10890
rect 1930 10650 2170 10890
rect 2260 10650 2500 10890
rect 2590 10650 2830 10890
rect 2920 10650 3160 10890
rect 3250 10650 3490 10890
rect 3580 10650 3820 10890
rect 3910 10650 4150 10890
rect 4240 10650 4480 10890
rect 4570 10650 4810 10890
rect 4900 10650 5140 10890
rect 5230 10650 5470 10890
rect 5560 10650 5800 10890
rect 5890 10650 6130 10890
rect 6220 10650 6460 10890
rect 6550 10650 6790 10890
rect 6880 10650 7120 10890
rect -4670 10320 -4430 10560
rect -4340 10320 -4100 10560
rect -4010 10320 -3770 10560
rect -3680 10320 -3440 10560
rect -3350 10320 -3110 10560
rect -3020 10320 -2780 10560
rect -2690 10320 -2450 10560
rect -2360 10320 -2120 10560
rect -2030 10320 -1790 10560
rect -1700 10320 -1460 10560
rect -1370 10320 -1130 10560
rect -1040 10320 -800 10560
rect -710 10320 -470 10560
rect -380 10320 -140 10560
rect -50 10320 190 10560
rect 280 10320 520 10560
rect 610 10320 850 10560
rect 940 10320 1180 10560
rect 1270 10320 1510 10560
rect 1600 10320 1840 10560
rect 1930 10320 2170 10560
rect 2260 10320 2500 10560
rect 2590 10320 2830 10560
rect 2920 10320 3160 10560
rect 3250 10320 3490 10560
rect 3580 10320 3820 10560
rect 3910 10320 4150 10560
rect 4240 10320 4480 10560
rect 4570 10320 4810 10560
rect 4900 10320 5140 10560
rect 5230 10320 5470 10560
rect 5560 10320 5800 10560
rect 5890 10320 6130 10560
rect 6220 10320 6460 10560
rect 6550 10320 6790 10560
rect 6880 10320 7120 10560
rect -4670 9990 -4430 10230
rect -4340 9990 -4100 10230
rect -4010 9990 -3770 10230
rect -3680 9990 -3440 10230
rect -3350 9990 -3110 10230
rect -3020 9990 -2780 10230
rect -2690 9990 -2450 10230
rect -2360 9990 -2120 10230
rect -2030 9990 -1790 10230
rect -1700 9990 -1460 10230
rect -1370 9990 -1130 10230
rect -1040 9990 -800 10230
rect -710 9990 -470 10230
rect -380 9990 -140 10230
rect -50 9990 190 10230
rect 280 9990 520 10230
rect 610 9990 850 10230
rect 940 9990 1180 10230
rect 1270 9990 1510 10230
rect 1600 9990 1840 10230
rect 1930 9990 2170 10230
rect 2260 9990 2500 10230
rect 2590 9990 2830 10230
rect 2920 9990 3160 10230
rect 3250 9990 3490 10230
rect 3580 9990 3820 10230
rect 3910 9990 4150 10230
rect 4240 9990 4480 10230
rect 4570 9990 4810 10230
rect 4900 9990 5140 10230
rect 5230 9990 5470 10230
rect 5560 9990 5800 10230
rect 5890 9990 6130 10230
rect 6220 9990 6460 10230
rect 6550 9990 6790 10230
rect 6880 9990 7120 10230
rect -4670 9660 -4430 9900
rect -4340 9660 -4100 9900
rect -4010 9660 -3770 9900
rect -3680 9660 -3440 9900
rect -3350 9660 -3110 9900
rect -3020 9660 -2780 9900
rect -2690 9660 -2450 9900
rect -2360 9660 -2120 9900
rect -2030 9660 -1790 9900
rect -1700 9660 -1460 9900
rect -1370 9660 -1130 9900
rect -1040 9660 -800 9900
rect -710 9660 -470 9900
rect -380 9660 -140 9900
rect -50 9660 190 9900
rect 280 9660 520 9900
rect 610 9660 850 9900
rect 940 9660 1180 9900
rect 1270 9660 1510 9900
rect 1600 9660 1840 9900
rect 1930 9660 2170 9900
rect 2260 9660 2500 9900
rect 2590 9660 2830 9900
rect 2920 9660 3160 9900
rect 3250 9660 3490 9900
rect 3580 9660 3820 9900
rect 3910 9660 4150 9900
rect 4240 9660 4480 9900
rect 4570 9660 4810 9900
rect 4900 9660 5140 9900
rect 5230 9660 5470 9900
rect 5560 9660 5800 9900
rect 5890 9660 6130 9900
rect 6220 9660 6460 9900
rect 6550 9660 6790 9900
rect 6880 9660 7120 9900
rect -4670 9330 -4430 9570
rect -4340 9330 -4100 9570
rect -4010 9330 -3770 9570
rect -3680 9330 -3440 9570
rect -3350 9330 -3110 9570
rect -3020 9330 -2780 9570
rect -2690 9330 -2450 9570
rect -2360 9330 -2120 9570
rect -2030 9330 -1790 9570
rect -1700 9330 -1460 9570
rect -1370 9330 -1130 9570
rect -1040 9330 -800 9570
rect -710 9330 -470 9570
rect -380 9330 -140 9570
rect -50 9330 190 9570
rect 280 9330 520 9570
rect 610 9330 850 9570
rect 940 9330 1180 9570
rect 1270 9330 1510 9570
rect 1600 9330 1840 9570
rect 1930 9330 2170 9570
rect 2260 9330 2500 9570
rect 2590 9330 2830 9570
rect 2920 9330 3160 9570
rect 3250 9330 3490 9570
rect 3580 9330 3820 9570
rect 3910 9330 4150 9570
rect 4240 9330 4480 9570
rect 4570 9330 4810 9570
rect 4900 9330 5140 9570
rect 5230 9330 5470 9570
rect 5560 9330 5800 9570
rect 5890 9330 6130 9570
rect 6220 9330 6460 9570
rect 6550 9330 6790 9570
rect 6880 9330 7120 9570
rect -4670 9000 -4430 9240
rect -4340 9000 -4100 9240
rect -4010 9000 -3770 9240
rect -3680 9000 -3440 9240
rect -3350 9000 -3110 9240
rect -3020 9000 -2780 9240
rect -2690 9000 -2450 9240
rect -2360 9000 -2120 9240
rect -2030 9000 -1790 9240
rect -1700 9000 -1460 9240
rect -1370 9000 -1130 9240
rect -1040 9000 -800 9240
rect -710 9000 -470 9240
rect -380 9000 -140 9240
rect -50 9000 190 9240
rect 280 9000 520 9240
rect 610 9000 850 9240
rect 940 9000 1180 9240
rect 1270 9000 1510 9240
rect 1600 9000 1840 9240
rect 1930 9000 2170 9240
rect 2260 9000 2500 9240
rect 2590 9000 2830 9240
rect 2920 9000 3160 9240
rect 3250 9000 3490 9240
rect 3580 9000 3820 9240
rect 3910 9000 4150 9240
rect 4240 9000 4480 9240
rect 4570 9000 4810 9240
rect 4900 9000 5140 9240
rect 5230 9000 5470 9240
rect 5560 9000 5800 9240
rect 5890 9000 6130 9240
rect 6220 9000 6460 9240
rect 6550 9000 6790 9240
rect 6880 9000 7120 9240
rect 7780 20550 8020 20790
rect 8110 20550 8350 20790
rect 8440 20550 8680 20790
rect 8770 20550 9010 20790
rect 9100 20550 9340 20790
rect 9430 20550 9670 20790
rect 9760 20550 10000 20790
rect 10090 20550 10330 20790
rect 10420 20550 10660 20790
rect 10750 20550 10990 20790
rect 11080 20550 11320 20790
rect 11410 20550 11650 20790
rect 11740 20550 11980 20790
rect 12070 20550 12310 20790
rect 12400 20550 12640 20790
rect 12730 20550 12970 20790
rect 13060 20550 13300 20790
rect 13390 20550 13630 20790
rect 13720 20550 13960 20790
rect 14050 20550 14290 20790
rect 14380 20550 14620 20790
rect 14710 20550 14950 20790
rect 15040 20550 15280 20790
rect 15370 20550 15610 20790
rect 15700 20550 15940 20790
rect 16030 20550 16270 20790
rect 16360 20550 16600 20790
rect 16690 20550 16930 20790
rect 17020 20550 17260 20790
rect 17350 20550 17590 20790
rect 17680 20550 17920 20790
rect 18010 20550 18250 20790
rect 18340 20550 18580 20790
rect 18670 20550 18910 20790
rect 19000 20550 19240 20790
rect 19330 20550 19570 20790
rect 7780 20220 8020 20460
rect 8110 20220 8350 20460
rect 8440 20220 8680 20460
rect 8770 20220 9010 20460
rect 9100 20220 9340 20460
rect 9430 20220 9670 20460
rect 9760 20220 10000 20460
rect 10090 20220 10330 20460
rect 10420 20220 10660 20460
rect 10750 20220 10990 20460
rect 11080 20220 11320 20460
rect 11410 20220 11650 20460
rect 11740 20220 11980 20460
rect 12070 20220 12310 20460
rect 12400 20220 12640 20460
rect 12730 20220 12970 20460
rect 13060 20220 13300 20460
rect 13390 20220 13630 20460
rect 13720 20220 13960 20460
rect 14050 20220 14290 20460
rect 14380 20220 14620 20460
rect 14710 20220 14950 20460
rect 15040 20220 15280 20460
rect 15370 20220 15610 20460
rect 15700 20220 15940 20460
rect 16030 20220 16270 20460
rect 16360 20220 16600 20460
rect 16690 20220 16930 20460
rect 17020 20220 17260 20460
rect 17350 20220 17590 20460
rect 17680 20220 17920 20460
rect 18010 20220 18250 20460
rect 18340 20220 18580 20460
rect 18670 20220 18910 20460
rect 19000 20220 19240 20460
rect 19330 20220 19570 20460
rect 7780 19890 8020 20130
rect 8110 19890 8350 20130
rect 8440 19890 8680 20130
rect 8770 19890 9010 20130
rect 9100 19890 9340 20130
rect 9430 19890 9670 20130
rect 9760 19890 10000 20130
rect 10090 19890 10330 20130
rect 10420 19890 10660 20130
rect 10750 19890 10990 20130
rect 11080 19890 11320 20130
rect 11410 19890 11650 20130
rect 11740 19890 11980 20130
rect 12070 19890 12310 20130
rect 12400 19890 12640 20130
rect 12730 19890 12970 20130
rect 13060 19890 13300 20130
rect 13390 19890 13630 20130
rect 13720 19890 13960 20130
rect 14050 19890 14290 20130
rect 14380 19890 14620 20130
rect 14710 19890 14950 20130
rect 15040 19890 15280 20130
rect 15370 19890 15610 20130
rect 15700 19890 15940 20130
rect 16030 19890 16270 20130
rect 16360 19890 16600 20130
rect 16690 19890 16930 20130
rect 17020 19890 17260 20130
rect 17350 19890 17590 20130
rect 17680 19890 17920 20130
rect 18010 19890 18250 20130
rect 18340 19890 18580 20130
rect 18670 19890 18910 20130
rect 19000 19890 19240 20130
rect 19330 19890 19570 20130
rect 7780 19560 8020 19800
rect 8110 19560 8350 19800
rect 8440 19560 8680 19800
rect 8770 19560 9010 19800
rect 9100 19560 9340 19800
rect 9430 19560 9670 19800
rect 9760 19560 10000 19800
rect 10090 19560 10330 19800
rect 10420 19560 10660 19800
rect 10750 19560 10990 19800
rect 11080 19560 11320 19800
rect 11410 19560 11650 19800
rect 11740 19560 11980 19800
rect 12070 19560 12310 19800
rect 12400 19560 12640 19800
rect 12730 19560 12970 19800
rect 13060 19560 13300 19800
rect 13390 19560 13630 19800
rect 13720 19560 13960 19800
rect 14050 19560 14290 19800
rect 14380 19560 14620 19800
rect 14710 19560 14950 19800
rect 15040 19560 15280 19800
rect 15370 19560 15610 19800
rect 15700 19560 15940 19800
rect 16030 19560 16270 19800
rect 16360 19560 16600 19800
rect 16690 19560 16930 19800
rect 17020 19560 17260 19800
rect 17350 19560 17590 19800
rect 17680 19560 17920 19800
rect 18010 19560 18250 19800
rect 18340 19560 18580 19800
rect 18670 19560 18910 19800
rect 19000 19560 19240 19800
rect 19330 19560 19570 19800
rect 7780 19230 8020 19470
rect 8110 19230 8350 19470
rect 8440 19230 8680 19470
rect 8770 19230 9010 19470
rect 9100 19230 9340 19470
rect 9430 19230 9670 19470
rect 9760 19230 10000 19470
rect 10090 19230 10330 19470
rect 10420 19230 10660 19470
rect 10750 19230 10990 19470
rect 11080 19230 11320 19470
rect 11410 19230 11650 19470
rect 11740 19230 11980 19470
rect 12070 19230 12310 19470
rect 12400 19230 12640 19470
rect 12730 19230 12970 19470
rect 13060 19230 13300 19470
rect 13390 19230 13630 19470
rect 13720 19230 13960 19470
rect 14050 19230 14290 19470
rect 14380 19230 14620 19470
rect 14710 19230 14950 19470
rect 15040 19230 15280 19470
rect 15370 19230 15610 19470
rect 15700 19230 15940 19470
rect 16030 19230 16270 19470
rect 16360 19230 16600 19470
rect 16690 19230 16930 19470
rect 17020 19230 17260 19470
rect 17350 19230 17590 19470
rect 17680 19230 17920 19470
rect 18010 19230 18250 19470
rect 18340 19230 18580 19470
rect 18670 19230 18910 19470
rect 19000 19230 19240 19470
rect 19330 19230 19570 19470
rect 7780 18900 8020 19140
rect 8110 18900 8350 19140
rect 8440 18900 8680 19140
rect 8770 18900 9010 19140
rect 9100 18900 9340 19140
rect 9430 18900 9670 19140
rect 9760 18900 10000 19140
rect 10090 18900 10330 19140
rect 10420 18900 10660 19140
rect 10750 18900 10990 19140
rect 11080 18900 11320 19140
rect 11410 18900 11650 19140
rect 11740 18900 11980 19140
rect 12070 18900 12310 19140
rect 12400 18900 12640 19140
rect 12730 18900 12970 19140
rect 13060 18900 13300 19140
rect 13390 18900 13630 19140
rect 13720 18900 13960 19140
rect 14050 18900 14290 19140
rect 14380 18900 14620 19140
rect 14710 18900 14950 19140
rect 15040 18900 15280 19140
rect 15370 18900 15610 19140
rect 15700 18900 15940 19140
rect 16030 18900 16270 19140
rect 16360 18900 16600 19140
rect 16690 18900 16930 19140
rect 17020 18900 17260 19140
rect 17350 18900 17590 19140
rect 17680 18900 17920 19140
rect 18010 18900 18250 19140
rect 18340 18900 18580 19140
rect 18670 18900 18910 19140
rect 19000 18900 19240 19140
rect 19330 18900 19570 19140
rect 7780 18570 8020 18810
rect 8110 18570 8350 18810
rect 8440 18570 8680 18810
rect 8770 18570 9010 18810
rect 9100 18570 9340 18810
rect 9430 18570 9670 18810
rect 9760 18570 10000 18810
rect 10090 18570 10330 18810
rect 10420 18570 10660 18810
rect 10750 18570 10990 18810
rect 11080 18570 11320 18810
rect 11410 18570 11650 18810
rect 11740 18570 11980 18810
rect 12070 18570 12310 18810
rect 12400 18570 12640 18810
rect 12730 18570 12970 18810
rect 13060 18570 13300 18810
rect 13390 18570 13630 18810
rect 13720 18570 13960 18810
rect 14050 18570 14290 18810
rect 14380 18570 14620 18810
rect 14710 18570 14950 18810
rect 15040 18570 15280 18810
rect 15370 18570 15610 18810
rect 15700 18570 15940 18810
rect 16030 18570 16270 18810
rect 16360 18570 16600 18810
rect 16690 18570 16930 18810
rect 17020 18570 17260 18810
rect 17350 18570 17590 18810
rect 17680 18570 17920 18810
rect 18010 18570 18250 18810
rect 18340 18570 18580 18810
rect 18670 18570 18910 18810
rect 19000 18570 19240 18810
rect 19330 18570 19570 18810
rect 7780 18240 8020 18480
rect 8110 18240 8350 18480
rect 8440 18240 8680 18480
rect 8770 18240 9010 18480
rect 9100 18240 9340 18480
rect 9430 18240 9670 18480
rect 9760 18240 10000 18480
rect 10090 18240 10330 18480
rect 10420 18240 10660 18480
rect 10750 18240 10990 18480
rect 11080 18240 11320 18480
rect 11410 18240 11650 18480
rect 11740 18240 11980 18480
rect 12070 18240 12310 18480
rect 12400 18240 12640 18480
rect 12730 18240 12970 18480
rect 13060 18240 13300 18480
rect 13390 18240 13630 18480
rect 13720 18240 13960 18480
rect 14050 18240 14290 18480
rect 14380 18240 14620 18480
rect 14710 18240 14950 18480
rect 15040 18240 15280 18480
rect 15370 18240 15610 18480
rect 15700 18240 15940 18480
rect 16030 18240 16270 18480
rect 16360 18240 16600 18480
rect 16690 18240 16930 18480
rect 17020 18240 17260 18480
rect 17350 18240 17590 18480
rect 17680 18240 17920 18480
rect 18010 18240 18250 18480
rect 18340 18240 18580 18480
rect 18670 18240 18910 18480
rect 19000 18240 19240 18480
rect 19330 18240 19570 18480
rect 7780 17910 8020 18150
rect 8110 17910 8350 18150
rect 8440 17910 8680 18150
rect 8770 17910 9010 18150
rect 9100 17910 9340 18150
rect 9430 17910 9670 18150
rect 9760 17910 10000 18150
rect 10090 17910 10330 18150
rect 10420 17910 10660 18150
rect 10750 17910 10990 18150
rect 11080 17910 11320 18150
rect 11410 17910 11650 18150
rect 11740 17910 11980 18150
rect 12070 17910 12310 18150
rect 12400 17910 12640 18150
rect 12730 17910 12970 18150
rect 13060 17910 13300 18150
rect 13390 17910 13630 18150
rect 13720 17910 13960 18150
rect 14050 17910 14290 18150
rect 14380 17910 14620 18150
rect 14710 17910 14950 18150
rect 15040 17910 15280 18150
rect 15370 17910 15610 18150
rect 15700 17910 15940 18150
rect 16030 17910 16270 18150
rect 16360 17910 16600 18150
rect 16690 17910 16930 18150
rect 17020 17910 17260 18150
rect 17350 17910 17590 18150
rect 17680 17910 17920 18150
rect 18010 17910 18250 18150
rect 18340 17910 18580 18150
rect 18670 17910 18910 18150
rect 19000 17910 19240 18150
rect 19330 17910 19570 18150
rect 7780 17580 8020 17820
rect 8110 17580 8350 17820
rect 8440 17580 8680 17820
rect 8770 17580 9010 17820
rect 9100 17580 9340 17820
rect 9430 17580 9670 17820
rect 9760 17580 10000 17820
rect 10090 17580 10330 17820
rect 10420 17580 10660 17820
rect 10750 17580 10990 17820
rect 11080 17580 11320 17820
rect 11410 17580 11650 17820
rect 11740 17580 11980 17820
rect 12070 17580 12310 17820
rect 12400 17580 12640 17820
rect 12730 17580 12970 17820
rect 13060 17580 13300 17820
rect 13390 17580 13630 17820
rect 13720 17580 13960 17820
rect 14050 17580 14290 17820
rect 14380 17580 14620 17820
rect 14710 17580 14950 17820
rect 15040 17580 15280 17820
rect 15370 17580 15610 17820
rect 15700 17580 15940 17820
rect 16030 17580 16270 17820
rect 16360 17580 16600 17820
rect 16690 17580 16930 17820
rect 17020 17580 17260 17820
rect 17350 17580 17590 17820
rect 17680 17580 17920 17820
rect 18010 17580 18250 17820
rect 18340 17580 18580 17820
rect 18670 17580 18910 17820
rect 19000 17580 19240 17820
rect 19330 17580 19570 17820
rect 7780 17250 8020 17490
rect 8110 17250 8350 17490
rect 8440 17250 8680 17490
rect 8770 17250 9010 17490
rect 9100 17250 9340 17490
rect 9430 17250 9670 17490
rect 9760 17250 10000 17490
rect 10090 17250 10330 17490
rect 10420 17250 10660 17490
rect 10750 17250 10990 17490
rect 11080 17250 11320 17490
rect 11410 17250 11650 17490
rect 11740 17250 11980 17490
rect 12070 17250 12310 17490
rect 12400 17250 12640 17490
rect 12730 17250 12970 17490
rect 13060 17250 13300 17490
rect 13390 17250 13630 17490
rect 13720 17250 13960 17490
rect 14050 17250 14290 17490
rect 14380 17250 14620 17490
rect 14710 17250 14950 17490
rect 15040 17250 15280 17490
rect 15370 17250 15610 17490
rect 15700 17250 15940 17490
rect 16030 17250 16270 17490
rect 16360 17250 16600 17490
rect 16690 17250 16930 17490
rect 17020 17250 17260 17490
rect 17350 17250 17590 17490
rect 17680 17250 17920 17490
rect 18010 17250 18250 17490
rect 18340 17250 18580 17490
rect 18670 17250 18910 17490
rect 19000 17250 19240 17490
rect 19330 17250 19570 17490
rect 7780 16920 8020 17160
rect 8110 16920 8350 17160
rect 8440 16920 8680 17160
rect 8770 16920 9010 17160
rect 9100 16920 9340 17160
rect 9430 16920 9670 17160
rect 9760 16920 10000 17160
rect 10090 16920 10330 17160
rect 10420 16920 10660 17160
rect 10750 16920 10990 17160
rect 11080 16920 11320 17160
rect 11410 16920 11650 17160
rect 11740 16920 11980 17160
rect 12070 16920 12310 17160
rect 12400 16920 12640 17160
rect 12730 16920 12970 17160
rect 13060 16920 13300 17160
rect 13390 16920 13630 17160
rect 13720 16920 13960 17160
rect 14050 16920 14290 17160
rect 14380 16920 14620 17160
rect 14710 16920 14950 17160
rect 15040 16920 15280 17160
rect 15370 16920 15610 17160
rect 15700 16920 15940 17160
rect 16030 16920 16270 17160
rect 16360 16920 16600 17160
rect 16690 16920 16930 17160
rect 17020 16920 17260 17160
rect 17350 16920 17590 17160
rect 17680 16920 17920 17160
rect 18010 16920 18250 17160
rect 18340 16920 18580 17160
rect 18670 16920 18910 17160
rect 19000 16920 19240 17160
rect 19330 16920 19570 17160
rect 7780 16590 8020 16830
rect 8110 16590 8350 16830
rect 8440 16590 8680 16830
rect 8770 16590 9010 16830
rect 9100 16590 9340 16830
rect 9430 16590 9670 16830
rect 9760 16590 10000 16830
rect 10090 16590 10330 16830
rect 10420 16590 10660 16830
rect 10750 16590 10990 16830
rect 11080 16590 11320 16830
rect 11410 16590 11650 16830
rect 11740 16590 11980 16830
rect 12070 16590 12310 16830
rect 12400 16590 12640 16830
rect 12730 16590 12970 16830
rect 13060 16590 13300 16830
rect 13390 16590 13630 16830
rect 13720 16590 13960 16830
rect 14050 16590 14290 16830
rect 14380 16590 14620 16830
rect 14710 16590 14950 16830
rect 15040 16590 15280 16830
rect 15370 16590 15610 16830
rect 15700 16590 15940 16830
rect 16030 16590 16270 16830
rect 16360 16590 16600 16830
rect 16690 16590 16930 16830
rect 17020 16590 17260 16830
rect 17350 16590 17590 16830
rect 17680 16590 17920 16830
rect 18010 16590 18250 16830
rect 18340 16590 18580 16830
rect 18670 16590 18910 16830
rect 19000 16590 19240 16830
rect 19330 16590 19570 16830
rect 7780 16260 8020 16500
rect 8110 16260 8350 16500
rect 8440 16260 8680 16500
rect 8770 16260 9010 16500
rect 9100 16260 9340 16500
rect 9430 16260 9670 16500
rect 9760 16260 10000 16500
rect 10090 16260 10330 16500
rect 10420 16260 10660 16500
rect 10750 16260 10990 16500
rect 11080 16260 11320 16500
rect 11410 16260 11650 16500
rect 11740 16260 11980 16500
rect 12070 16260 12310 16500
rect 12400 16260 12640 16500
rect 12730 16260 12970 16500
rect 13060 16260 13300 16500
rect 13390 16260 13630 16500
rect 13720 16260 13960 16500
rect 14050 16260 14290 16500
rect 14380 16260 14620 16500
rect 14710 16260 14950 16500
rect 15040 16260 15280 16500
rect 15370 16260 15610 16500
rect 15700 16260 15940 16500
rect 16030 16260 16270 16500
rect 16360 16260 16600 16500
rect 16690 16260 16930 16500
rect 17020 16260 17260 16500
rect 17350 16260 17590 16500
rect 17680 16260 17920 16500
rect 18010 16260 18250 16500
rect 18340 16260 18580 16500
rect 18670 16260 18910 16500
rect 19000 16260 19240 16500
rect 19330 16260 19570 16500
rect 7780 15930 8020 16170
rect 8110 15930 8350 16170
rect 8440 15930 8680 16170
rect 8770 15930 9010 16170
rect 9100 15930 9340 16170
rect 9430 15930 9670 16170
rect 9760 15930 10000 16170
rect 10090 15930 10330 16170
rect 10420 15930 10660 16170
rect 10750 15930 10990 16170
rect 11080 15930 11320 16170
rect 11410 15930 11650 16170
rect 11740 15930 11980 16170
rect 12070 15930 12310 16170
rect 12400 15930 12640 16170
rect 12730 15930 12970 16170
rect 13060 15930 13300 16170
rect 13390 15930 13630 16170
rect 13720 15930 13960 16170
rect 14050 15930 14290 16170
rect 14380 15930 14620 16170
rect 14710 15930 14950 16170
rect 15040 15930 15280 16170
rect 15370 15930 15610 16170
rect 15700 15930 15940 16170
rect 16030 15930 16270 16170
rect 16360 15930 16600 16170
rect 16690 15930 16930 16170
rect 17020 15930 17260 16170
rect 17350 15930 17590 16170
rect 17680 15930 17920 16170
rect 18010 15930 18250 16170
rect 18340 15930 18580 16170
rect 18670 15930 18910 16170
rect 19000 15930 19240 16170
rect 19330 15930 19570 16170
rect 7780 15600 8020 15840
rect 8110 15600 8350 15840
rect 8440 15600 8680 15840
rect 8770 15600 9010 15840
rect 9100 15600 9340 15840
rect 9430 15600 9670 15840
rect 9760 15600 10000 15840
rect 10090 15600 10330 15840
rect 10420 15600 10660 15840
rect 10750 15600 10990 15840
rect 11080 15600 11320 15840
rect 11410 15600 11650 15840
rect 11740 15600 11980 15840
rect 12070 15600 12310 15840
rect 12400 15600 12640 15840
rect 12730 15600 12970 15840
rect 13060 15600 13300 15840
rect 13390 15600 13630 15840
rect 13720 15600 13960 15840
rect 14050 15600 14290 15840
rect 14380 15600 14620 15840
rect 14710 15600 14950 15840
rect 15040 15600 15280 15840
rect 15370 15600 15610 15840
rect 15700 15600 15940 15840
rect 16030 15600 16270 15840
rect 16360 15600 16600 15840
rect 16690 15600 16930 15840
rect 17020 15600 17260 15840
rect 17350 15600 17590 15840
rect 17680 15600 17920 15840
rect 18010 15600 18250 15840
rect 18340 15600 18580 15840
rect 18670 15600 18910 15840
rect 19000 15600 19240 15840
rect 19330 15600 19570 15840
rect 7780 15270 8020 15510
rect 8110 15270 8350 15510
rect 8440 15270 8680 15510
rect 8770 15270 9010 15510
rect 9100 15270 9340 15510
rect 9430 15270 9670 15510
rect 9760 15270 10000 15510
rect 10090 15270 10330 15510
rect 10420 15270 10660 15510
rect 10750 15270 10990 15510
rect 11080 15270 11320 15510
rect 11410 15270 11650 15510
rect 11740 15270 11980 15510
rect 12070 15270 12310 15510
rect 12400 15270 12640 15510
rect 12730 15270 12970 15510
rect 13060 15270 13300 15510
rect 13390 15270 13630 15510
rect 13720 15270 13960 15510
rect 14050 15270 14290 15510
rect 14380 15270 14620 15510
rect 14710 15270 14950 15510
rect 15040 15270 15280 15510
rect 15370 15270 15610 15510
rect 15700 15270 15940 15510
rect 16030 15270 16270 15510
rect 16360 15270 16600 15510
rect 16690 15270 16930 15510
rect 17020 15270 17260 15510
rect 17350 15270 17590 15510
rect 17680 15270 17920 15510
rect 18010 15270 18250 15510
rect 18340 15270 18580 15510
rect 18670 15270 18910 15510
rect 19000 15270 19240 15510
rect 19330 15270 19570 15510
rect 7780 14940 8020 15180
rect 8110 14940 8350 15180
rect 8440 14940 8680 15180
rect 8770 14940 9010 15180
rect 9100 14940 9340 15180
rect 9430 14940 9670 15180
rect 9760 14940 10000 15180
rect 10090 14940 10330 15180
rect 10420 14940 10660 15180
rect 10750 14940 10990 15180
rect 11080 14940 11320 15180
rect 11410 14940 11650 15180
rect 11740 14940 11980 15180
rect 12070 14940 12310 15180
rect 12400 14940 12640 15180
rect 12730 14940 12970 15180
rect 13060 14940 13300 15180
rect 13390 14940 13630 15180
rect 13720 14940 13960 15180
rect 14050 14940 14290 15180
rect 14380 14940 14620 15180
rect 14710 14940 14950 15180
rect 15040 14940 15280 15180
rect 15370 14940 15610 15180
rect 15700 14940 15940 15180
rect 16030 14940 16270 15180
rect 16360 14940 16600 15180
rect 16690 14940 16930 15180
rect 17020 14940 17260 15180
rect 17350 14940 17590 15180
rect 17680 14940 17920 15180
rect 18010 14940 18250 15180
rect 18340 14940 18580 15180
rect 18670 14940 18910 15180
rect 19000 14940 19240 15180
rect 19330 14940 19570 15180
rect 7780 14610 8020 14850
rect 8110 14610 8350 14850
rect 8440 14610 8680 14850
rect 8770 14610 9010 14850
rect 9100 14610 9340 14850
rect 9430 14610 9670 14850
rect 9760 14610 10000 14850
rect 10090 14610 10330 14850
rect 10420 14610 10660 14850
rect 10750 14610 10990 14850
rect 11080 14610 11320 14850
rect 11410 14610 11650 14850
rect 11740 14610 11980 14850
rect 12070 14610 12310 14850
rect 12400 14610 12640 14850
rect 12730 14610 12970 14850
rect 13060 14610 13300 14850
rect 13390 14610 13630 14850
rect 13720 14610 13960 14850
rect 14050 14610 14290 14850
rect 14380 14610 14620 14850
rect 14710 14610 14950 14850
rect 15040 14610 15280 14850
rect 15370 14610 15610 14850
rect 15700 14610 15940 14850
rect 16030 14610 16270 14850
rect 16360 14610 16600 14850
rect 16690 14610 16930 14850
rect 17020 14610 17260 14850
rect 17350 14610 17590 14850
rect 17680 14610 17920 14850
rect 18010 14610 18250 14850
rect 18340 14610 18580 14850
rect 18670 14610 18910 14850
rect 19000 14610 19240 14850
rect 19330 14610 19570 14850
rect 7780 14280 8020 14520
rect 8110 14280 8350 14520
rect 8440 14280 8680 14520
rect 8770 14280 9010 14520
rect 9100 14280 9340 14520
rect 9430 14280 9670 14520
rect 9760 14280 10000 14520
rect 10090 14280 10330 14520
rect 10420 14280 10660 14520
rect 10750 14280 10990 14520
rect 11080 14280 11320 14520
rect 11410 14280 11650 14520
rect 11740 14280 11980 14520
rect 12070 14280 12310 14520
rect 12400 14280 12640 14520
rect 12730 14280 12970 14520
rect 13060 14280 13300 14520
rect 13390 14280 13630 14520
rect 13720 14280 13960 14520
rect 14050 14280 14290 14520
rect 14380 14280 14620 14520
rect 14710 14280 14950 14520
rect 15040 14280 15280 14520
rect 15370 14280 15610 14520
rect 15700 14280 15940 14520
rect 16030 14280 16270 14520
rect 16360 14280 16600 14520
rect 16690 14280 16930 14520
rect 17020 14280 17260 14520
rect 17350 14280 17590 14520
rect 17680 14280 17920 14520
rect 18010 14280 18250 14520
rect 18340 14280 18580 14520
rect 18670 14280 18910 14520
rect 19000 14280 19240 14520
rect 19330 14280 19570 14520
rect 7780 13950 8020 14190
rect 8110 13950 8350 14190
rect 8440 13950 8680 14190
rect 8770 13950 9010 14190
rect 9100 13950 9340 14190
rect 9430 13950 9670 14190
rect 9760 13950 10000 14190
rect 10090 13950 10330 14190
rect 10420 13950 10660 14190
rect 10750 13950 10990 14190
rect 11080 13950 11320 14190
rect 11410 13950 11650 14190
rect 11740 13950 11980 14190
rect 12070 13950 12310 14190
rect 12400 13950 12640 14190
rect 12730 13950 12970 14190
rect 13060 13950 13300 14190
rect 13390 13950 13630 14190
rect 13720 13950 13960 14190
rect 14050 13950 14290 14190
rect 14380 13950 14620 14190
rect 14710 13950 14950 14190
rect 15040 13950 15280 14190
rect 15370 13950 15610 14190
rect 15700 13950 15940 14190
rect 16030 13950 16270 14190
rect 16360 13950 16600 14190
rect 16690 13950 16930 14190
rect 17020 13950 17260 14190
rect 17350 13950 17590 14190
rect 17680 13950 17920 14190
rect 18010 13950 18250 14190
rect 18340 13950 18580 14190
rect 18670 13950 18910 14190
rect 19000 13950 19240 14190
rect 19330 13950 19570 14190
rect 7780 13620 8020 13860
rect 8110 13620 8350 13860
rect 8440 13620 8680 13860
rect 8770 13620 9010 13860
rect 9100 13620 9340 13860
rect 9430 13620 9670 13860
rect 9760 13620 10000 13860
rect 10090 13620 10330 13860
rect 10420 13620 10660 13860
rect 10750 13620 10990 13860
rect 11080 13620 11320 13860
rect 11410 13620 11650 13860
rect 11740 13620 11980 13860
rect 12070 13620 12310 13860
rect 12400 13620 12640 13860
rect 12730 13620 12970 13860
rect 13060 13620 13300 13860
rect 13390 13620 13630 13860
rect 13720 13620 13960 13860
rect 14050 13620 14290 13860
rect 14380 13620 14620 13860
rect 14710 13620 14950 13860
rect 15040 13620 15280 13860
rect 15370 13620 15610 13860
rect 15700 13620 15940 13860
rect 16030 13620 16270 13860
rect 16360 13620 16600 13860
rect 16690 13620 16930 13860
rect 17020 13620 17260 13860
rect 17350 13620 17590 13860
rect 17680 13620 17920 13860
rect 18010 13620 18250 13860
rect 18340 13620 18580 13860
rect 18670 13620 18910 13860
rect 19000 13620 19240 13860
rect 19330 13620 19570 13860
rect 7780 13290 8020 13530
rect 8110 13290 8350 13530
rect 8440 13290 8680 13530
rect 8770 13290 9010 13530
rect 9100 13290 9340 13530
rect 9430 13290 9670 13530
rect 9760 13290 10000 13530
rect 10090 13290 10330 13530
rect 10420 13290 10660 13530
rect 10750 13290 10990 13530
rect 11080 13290 11320 13530
rect 11410 13290 11650 13530
rect 11740 13290 11980 13530
rect 12070 13290 12310 13530
rect 12400 13290 12640 13530
rect 12730 13290 12970 13530
rect 13060 13290 13300 13530
rect 13390 13290 13630 13530
rect 13720 13290 13960 13530
rect 14050 13290 14290 13530
rect 14380 13290 14620 13530
rect 14710 13290 14950 13530
rect 15040 13290 15280 13530
rect 15370 13290 15610 13530
rect 15700 13290 15940 13530
rect 16030 13290 16270 13530
rect 16360 13290 16600 13530
rect 16690 13290 16930 13530
rect 17020 13290 17260 13530
rect 17350 13290 17590 13530
rect 17680 13290 17920 13530
rect 18010 13290 18250 13530
rect 18340 13290 18580 13530
rect 18670 13290 18910 13530
rect 19000 13290 19240 13530
rect 19330 13290 19570 13530
rect 7780 12960 8020 13200
rect 8110 12960 8350 13200
rect 8440 12960 8680 13200
rect 8770 12960 9010 13200
rect 9100 12960 9340 13200
rect 9430 12960 9670 13200
rect 9760 12960 10000 13200
rect 10090 12960 10330 13200
rect 10420 12960 10660 13200
rect 10750 12960 10990 13200
rect 11080 12960 11320 13200
rect 11410 12960 11650 13200
rect 11740 12960 11980 13200
rect 12070 12960 12310 13200
rect 12400 12960 12640 13200
rect 12730 12960 12970 13200
rect 13060 12960 13300 13200
rect 13390 12960 13630 13200
rect 13720 12960 13960 13200
rect 14050 12960 14290 13200
rect 14380 12960 14620 13200
rect 14710 12960 14950 13200
rect 15040 12960 15280 13200
rect 15370 12960 15610 13200
rect 15700 12960 15940 13200
rect 16030 12960 16270 13200
rect 16360 12960 16600 13200
rect 16690 12960 16930 13200
rect 17020 12960 17260 13200
rect 17350 12960 17590 13200
rect 17680 12960 17920 13200
rect 18010 12960 18250 13200
rect 18340 12960 18580 13200
rect 18670 12960 18910 13200
rect 19000 12960 19240 13200
rect 19330 12960 19570 13200
rect 7780 12630 8020 12870
rect 8110 12630 8350 12870
rect 8440 12630 8680 12870
rect 8770 12630 9010 12870
rect 9100 12630 9340 12870
rect 9430 12630 9670 12870
rect 9760 12630 10000 12870
rect 10090 12630 10330 12870
rect 10420 12630 10660 12870
rect 10750 12630 10990 12870
rect 11080 12630 11320 12870
rect 11410 12630 11650 12870
rect 11740 12630 11980 12870
rect 12070 12630 12310 12870
rect 12400 12630 12640 12870
rect 12730 12630 12970 12870
rect 13060 12630 13300 12870
rect 13390 12630 13630 12870
rect 13720 12630 13960 12870
rect 14050 12630 14290 12870
rect 14380 12630 14620 12870
rect 14710 12630 14950 12870
rect 15040 12630 15280 12870
rect 15370 12630 15610 12870
rect 15700 12630 15940 12870
rect 16030 12630 16270 12870
rect 16360 12630 16600 12870
rect 16690 12630 16930 12870
rect 17020 12630 17260 12870
rect 17350 12630 17590 12870
rect 17680 12630 17920 12870
rect 18010 12630 18250 12870
rect 18340 12630 18580 12870
rect 18670 12630 18910 12870
rect 19000 12630 19240 12870
rect 19330 12630 19570 12870
rect 7780 12300 8020 12540
rect 8110 12300 8350 12540
rect 8440 12300 8680 12540
rect 8770 12300 9010 12540
rect 9100 12300 9340 12540
rect 9430 12300 9670 12540
rect 9760 12300 10000 12540
rect 10090 12300 10330 12540
rect 10420 12300 10660 12540
rect 10750 12300 10990 12540
rect 11080 12300 11320 12540
rect 11410 12300 11650 12540
rect 11740 12300 11980 12540
rect 12070 12300 12310 12540
rect 12400 12300 12640 12540
rect 12730 12300 12970 12540
rect 13060 12300 13300 12540
rect 13390 12300 13630 12540
rect 13720 12300 13960 12540
rect 14050 12300 14290 12540
rect 14380 12300 14620 12540
rect 14710 12300 14950 12540
rect 15040 12300 15280 12540
rect 15370 12300 15610 12540
rect 15700 12300 15940 12540
rect 16030 12300 16270 12540
rect 16360 12300 16600 12540
rect 16690 12300 16930 12540
rect 17020 12300 17260 12540
rect 17350 12300 17590 12540
rect 17680 12300 17920 12540
rect 18010 12300 18250 12540
rect 18340 12300 18580 12540
rect 18670 12300 18910 12540
rect 19000 12300 19240 12540
rect 19330 12300 19570 12540
rect 7780 11970 8020 12210
rect 8110 11970 8350 12210
rect 8440 11970 8680 12210
rect 8770 11970 9010 12210
rect 9100 11970 9340 12210
rect 9430 11970 9670 12210
rect 9760 11970 10000 12210
rect 10090 11970 10330 12210
rect 10420 11970 10660 12210
rect 10750 11970 10990 12210
rect 11080 11970 11320 12210
rect 11410 11970 11650 12210
rect 11740 11970 11980 12210
rect 12070 11970 12310 12210
rect 12400 11970 12640 12210
rect 12730 11970 12970 12210
rect 13060 11970 13300 12210
rect 13390 11970 13630 12210
rect 13720 11970 13960 12210
rect 14050 11970 14290 12210
rect 14380 11970 14620 12210
rect 14710 11970 14950 12210
rect 15040 11970 15280 12210
rect 15370 11970 15610 12210
rect 15700 11970 15940 12210
rect 16030 11970 16270 12210
rect 16360 11970 16600 12210
rect 16690 11970 16930 12210
rect 17020 11970 17260 12210
rect 17350 11970 17590 12210
rect 17680 11970 17920 12210
rect 18010 11970 18250 12210
rect 18340 11970 18580 12210
rect 18670 11970 18910 12210
rect 19000 11970 19240 12210
rect 19330 11970 19570 12210
rect 7780 11640 8020 11880
rect 8110 11640 8350 11880
rect 8440 11640 8680 11880
rect 8770 11640 9010 11880
rect 9100 11640 9340 11880
rect 9430 11640 9670 11880
rect 9760 11640 10000 11880
rect 10090 11640 10330 11880
rect 10420 11640 10660 11880
rect 10750 11640 10990 11880
rect 11080 11640 11320 11880
rect 11410 11640 11650 11880
rect 11740 11640 11980 11880
rect 12070 11640 12310 11880
rect 12400 11640 12640 11880
rect 12730 11640 12970 11880
rect 13060 11640 13300 11880
rect 13390 11640 13630 11880
rect 13720 11640 13960 11880
rect 14050 11640 14290 11880
rect 14380 11640 14620 11880
rect 14710 11640 14950 11880
rect 15040 11640 15280 11880
rect 15370 11640 15610 11880
rect 15700 11640 15940 11880
rect 16030 11640 16270 11880
rect 16360 11640 16600 11880
rect 16690 11640 16930 11880
rect 17020 11640 17260 11880
rect 17350 11640 17590 11880
rect 17680 11640 17920 11880
rect 18010 11640 18250 11880
rect 18340 11640 18580 11880
rect 18670 11640 18910 11880
rect 19000 11640 19240 11880
rect 19330 11640 19570 11880
rect 7780 11310 8020 11550
rect 8110 11310 8350 11550
rect 8440 11310 8680 11550
rect 8770 11310 9010 11550
rect 9100 11310 9340 11550
rect 9430 11310 9670 11550
rect 9760 11310 10000 11550
rect 10090 11310 10330 11550
rect 10420 11310 10660 11550
rect 10750 11310 10990 11550
rect 11080 11310 11320 11550
rect 11410 11310 11650 11550
rect 11740 11310 11980 11550
rect 12070 11310 12310 11550
rect 12400 11310 12640 11550
rect 12730 11310 12970 11550
rect 13060 11310 13300 11550
rect 13390 11310 13630 11550
rect 13720 11310 13960 11550
rect 14050 11310 14290 11550
rect 14380 11310 14620 11550
rect 14710 11310 14950 11550
rect 15040 11310 15280 11550
rect 15370 11310 15610 11550
rect 15700 11310 15940 11550
rect 16030 11310 16270 11550
rect 16360 11310 16600 11550
rect 16690 11310 16930 11550
rect 17020 11310 17260 11550
rect 17350 11310 17590 11550
rect 17680 11310 17920 11550
rect 18010 11310 18250 11550
rect 18340 11310 18580 11550
rect 18670 11310 18910 11550
rect 19000 11310 19240 11550
rect 19330 11310 19570 11550
rect 7780 10980 8020 11220
rect 8110 10980 8350 11220
rect 8440 10980 8680 11220
rect 8770 10980 9010 11220
rect 9100 10980 9340 11220
rect 9430 10980 9670 11220
rect 9760 10980 10000 11220
rect 10090 10980 10330 11220
rect 10420 10980 10660 11220
rect 10750 10980 10990 11220
rect 11080 10980 11320 11220
rect 11410 10980 11650 11220
rect 11740 10980 11980 11220
rect 12070 10980 12310 11220
rect 12400 10980 12640 11220
rect 12730 10980 12970 11220
rect 13060 10980 13300 11220
rect 13390 10980 13630 11220
rect 13720 10980 13960 11220
rect 14050 10980 14290 11220
rect 14380 10980 14620 11220
rect 14710 10980 14950 11220
rect 15040 10980 15280 11220
rect 15370 10980 15610 11220
rect 15700 10980 15940 11220
rect 16030 10980 16270 11220
rect 16360 10980 16600 11220
rect 16690 10980 16930 11220
rect 17020 10980 17260 11220
rect 17350 10980 17590 11220
rect 17680 10980 17920 11220
rect 18010 10980 18250 11220
rect 18340 10980 18580 11220
rect 18670 10980 18910 11220
rect 19000 10980 19240 11220
rect 19330 10980 19570 11220
rect 7780 10650 8020 10890
rect 8110 10650 8350 10890
rect 8440 10650 8680 10890
rect 8770 10650 9010 10890
rect 9100 10650 9340 10890
rect 9430 10650 9670 10890
rect 9760 10650 10000 10890
rect 10090 10650 10330 10890
rect 10420 10650 10660 10890
rect 10750 10650 10990 10890
rect 11080 10650 11320 10890
rect 11410 10650 11650 10890
rect 11740 10650 11980 10890
rect 12070 10650 12310 10890
rect 12400 10650 12640 10890
rect 12730 10650 12970 10890
rect 13060 10650 13300 10890
rect 13390 10650 13630 10890
rect 13720 10650 13960 10890
rect 14050 10650 14290 10890
rect 14380 10650 14620 10890
rect 14710 10650 14950 10890
rect 15040 10650 15280 10890
rect 15370 10650 15610 10890
rect 15700 10650 15940 10890
rect 16030 10650 16270 10890
rect 16360 10650 16600 10890
rect 16690 10650 16930 10890
rect 17020 10650 17260 10890
rect 17350 10650 17590 10890
rect 17680 10650 17920 10890
rect 18010 10650 18250 10890
rect 18340 10650 18580 10890
rect 18670 10650 18910 10890
rect 19000 10650 19240 10890
rect 19330 10650 19570 10890
rect 7780 10320 8020 10560
rect 8110 10320 8350 10560
rect 8440 10320 8680 10560
rect 8770 10320 9010 10560
rect 9100 10320 9340 10560
rect 9430 10320 9670 10560
rect 9760 10320 10000 10560
rect 10090 10320 10330 10560
rect 10420 10320 10660 10560
rect 10750 10320 10990 10560
rect 11080 10320 11320 10560
rect 11410 10320 11650 10560
rect 11740 10320 11980 10560
rect 12070 10320 12310 10560
rect 12400 10320 12640 10560
rect 12730 10320 12970 10560
rect 13060 10320 13300 10560
rect 13390 10320 13630 10560
rect 13720 10320 13960 10560
rect 14050 10320 14290 10560
rect 14380 10320 14620 10560
rect 14710 10320 14950 10560
rect 15040 10320 15280 10560
rect 15370 10320 15610 10560
rect 15700 10320 15940 10560
rect 16030 10320 16270 10560
rect 16360 10320 16600 10560
rect 16690 10320 16930 10560
rect 17020 10320 17260 10560
rect 17350 10320 17590 10560
rect 17680 10320 17920 10560
rect 18010 10320 18250 10560
rect 18340 10320 18580 10560
rect 18670 10320 18910 10560
rect 19000 10320 19240 10560
rect 19330 10320 19570 10560
rect 7780 9990 8020 10230
rect 8110 9990 8350 10230
rect 8440 9990 8680 10230
rect 8770 9990 9010 10230
rect 9100 9990 9340 10230
rect 9430 9990 9670 10230
rect 9760 9990 10000 10230
rect 10090 9990 10330 10230
rect 10420 9990 10660 10230
rect 10750 9990 10990 10230
rect 11080 9990 11320 10230
rect 11410 9990 11650 10230
rect 11740 9990 11980 10230
rect 12070 9990 12310 10230
rect 12400 9990 12640 10230
rect 12730 9990 12970 10230
rect 13060 9990 13300 10230
rect 13390 9990 13630 10230
rect 13720 9990 13960 10230
rect 14050 9990 14290 10230
rect 14380 9990 14620 10230
rect 14710 9990 14950 10230
rect 15040 9990 15280 10230
rect 15370 9990 15610 10230
rect 15700 9990 15940 10230
rect 16030 9990 16270 10230
rect 16360 9990 16600 10230
rect 16690 9990 16930 10230
rect 17020 9990 17260 10230
rect 17350 9990 17590 10230
rect 17680 9990 17920 10230
rect 18010 9990 18250 10230
rect 18340 9990 18580 10230
rect 18670 9990 18910 10230
rect 19000 9990 19240 10230
rect 19330 9990 19570 10230
rect 7780 9660 8020 9900
rect 8110 9660 8350 9900
rect 8440 9660 8680 9900
rect 8770 9660 9010 9900
rect 9100 9660 9340 9900
rect 9430 9660 9670 9900
rect 9760 9660 10000 9900
rect 10090 9660 10330 9900
rect 10420 9660 10660 9900
rect 10750 9660 10990 9900
rect 11080 9660 11320 9900
rect 11410 9660 11650 9900
rect 11740 9660 11980 9900
rect 12070 9660 12310 9900
rect 12400 9660 12640 9900
rect 12730 9660 12970 9900
rect 13060 9660 13300 9900
rect 13390 9660 13630 9900
rect 13720 9660 13960 9900
rect 14050 9660 14290 9900
rect 14380 9660 14620 9900
rect 14710 9660 14950 9900
rect 15040 9660 15280 9900
rect 15370 9660 15610 9900
rect 15700 9660 15940 9900
rect 16030 9660 16270 9900
rect 16360 9660 16600 9900
rect 16690 9660 16930 9900
rect 17020 9660 17260 9900
rect 17350 9660 17590 9900
rect 17680 9660 17920 9900
rect 18010 9660 18250 9900
rect 18340 9660 18580 9900
rect 18670 9660 18910 9900
rect 19000 9660 19240 9900
rect 19330 9660 19570 9900
rect 7780 9330 8020 9570
rect 8110 9330 8350 9570
rect 8440 9330 8680 9570
rect 8770 9330 9010 9570
rect 9100 9330 9340 9570
rect 9430 9330 9670 9570
rect 9760 9330 10000 9570
rect 10090 9330 10330 9570
rect 10420 9330 10660 9570
rect 10750 9330 10990 9570
rect 11080 9330 11320 9570
rect 11410 9330 11650 9570
rect 11740 9330 11980 9570
rect 12070 9330 12310 9570
rect 12400 9330 12640 9570
rect 12730 9330 12970 9570
rect 13060 9330 13300 9570
rect 13390 9330 13630 9570
rect 13720 9330 13960 9570
rect 14050 9330 14290 9570
rect 14380 9330 14620 9570
rect 14710 9330 14950 9570
rect 15040 9330 15280 9570
rect 15370 9330 15610 9570
rect 15700 9330 15940 9570
rect 16030 9330 16270 9570
rect 16360 9330 16600 9570
rect 16690 9330 16930 9570
rect 17020 9330 17260 9570
rect 17350 9330 17590 9570
rect 17680 9330 17920 9570
rect 18010 9330 18250 9570
rect 18340 9330 18580 9570
rect 18670 9330 18910 9570
rect 19000 9330 19240 9570
rect 19330 9330 19570 9570
rect 7780 9000 8020 9240
rect 8110 9000 8350 9240
rect 8440 9000 8680 9240
rect 8770 9000 9010 9240
rect 9100 9000 9340 9240
rect 9430 9000 9670 9240
rect 9760 9000 10000 9240
rect 10090 9000 10330 9240
rect 10420 9000 10660 9240
rect 10750 9000 10990 9240
rect 11080 9000 11320 9240
rect 11410 9000 11650 9240
rect 11740 9000 11980 9240
rect 12070 9000 12310 9240
rect 12400 9000 12640 9240
rect 12730 9000 12970 9240
rect 13060 9000 13300 9240
rect 13390 9000 13630 9240
rect 13720 9000 13960 9240
rect 14050 9000 14290 9240
rect 14380 9000 14620 9240
rect 14710 9000 14950 9240
rect 15040 9000 15280 9240
rect 15370 9000 15610 9240
rect 15700 9000 15940 9240
rect 16030 9000 16270 9240
rect 16360 9000 16600 9240
rect 16690 9000 16930 9240
rect 17020 9000 17260 9240
rect 17350 9000 17590 9240
rect 17680 9000 17920 9240
rect 18010 9000 18250 9240
rect 18340 9000 18580 9240
rect 18670 9000 18910 9240
rect 19000 9000 19240 9240
rect 19330 9000 19570 9240
rect 28780 7590 29020 7830
rect 29110 7590 29350 7830
rect 29440 7590 29680 7830
rect 29770 7590 30010 7830
rect 30100 7590 30340 7830
rect 30430 7590 30670 7830
rect 30760 7590 31000 7830
rect 31090 7590 31330 7830
rect 31420 7590 31660 7830
rect 31750 7590 31990 7830
rect 32080 7590 32320 7830
rect 32410 7590 32650 7830
rect 32740 7590 32980 7830
rect 33070 7590 33310 7830
rect 33400 7590 33640 7830
rect 33730 7590 33970 7830
rect 34060 7590 34300 7830
rect 34390 7590 34630 7830
rect 34720 7590 34960 7830
rect 35050 7590 35290 7830
rect 28780 7260 29020 7500
rect 29110 7260 29350 7500
rect 29440 7260 29680 7500
rect 29770 7260 30010 7500
rect 30100 7260 30340 7500
rect 30430 7260 30670 7500
rect 30760 7260 31000 7500
rect 31090 7260 31330 7500
rect 31420 7260 31660 7500
rect 31750 7260 31990 7500
rect 32080 7260 32320 7500
rect 32410 7260 32650 7500
rect 32740 7260 32980 7500
rect 33070 7260 33310 7500
rect 33400 7260 33640 7500
rect 33730 7260 33970 7500
rect 34060 7260 34300 7500
rect 34390 7260 34630 7500
rect 34720 7260 34960 7500
rect 35050 7260 35290 7500
rect 28780 6930 29020 7170
rect 29110 6930 29350 7170
rect 29440 6930 29680 7170
rect 29770 6930 30010 7170
rect 30100 6930 30340 7170
rect 30430 6930 30670 7170
rect 30760 6930 31000 7170
rect 31090 6930 31330 7170
rect 31420 6930 31660 7170
rect 31750 6930 31990 7170
rect 32080 6930 32320 7170
rect 32410 6930 32650 7170
rect 32740 6930 32980 7170
rect 33070 6930 33310 7170
rect 33400 6930 33640 7170
rect 33730 6930 33970 7170
rect 34060 6930 34300 7170
rect 34390 6930 34630 7170
rect 34720 6930 34960 7170
rect 35050 6930 35290 7170
rect 28780 6600 29020 6840
rect 29110 6600 29350 6840
rect 29440 6600 29680 6840
rect 29770 6600 30010 6840
rect 30100 6600 30340 6840
rect 30430 6600 30670 6840
rect 30760 6600 31000 6840
rect 31090 6600 31330 6840
rect 31420 6600 31660 6840
rect 31750 6600 31990 6840
rect 32080 6600 32320 6840
rect 32410 6600 32650 6840
rect 32740 6600 32980 6840
rect 33070 6600 33310 6840
rect 33400 6600 33640 6840
rect 33730 6600 33970 6840
rect 34060 6600 34300 6840
rect 34390 6600 34630 6840
rect 34720 6600 34960 6840
rect 35050 6600 35290 6840
rect 28780 6270 29020 6510
rect 29110 6270 29350 6510
rect 29440 6270 29680 6510
rect 29770 6270 30010 6510
rect 30100 6270 30340 6510
rect 30430 6270 30670 6510
rect 30760 6270 31000 6510
rect 31090 6270 31330 6510
rect 31420 6270 31660 6510
rect 31750 6270 31990 6510
rect 32080 6270 32320 6510
rect 32410 6270 32650 6510
rect 32740 6270 32980 6510
rect 33070 6270 33310 6510
rect 33400 6270 33640 6510
rect 33730 6270 33970 6510
rect 34060 6270 34300 6510
rect 34390 6270 34630 6510
rect 34720 6270 34960 6510
rect 35050 6270 35290 6510
rect 28780 5940 29020 6180
rect 29110 5940 29350 6180
rect 29440 5940 29680 6180
rect 29770 5940 30010 6180
rect 30100 5940 30340 6180
rect 30430 5940 30670 6180
rect 30760 5940 31000 6180
rect 31090 5940 31330 6180
rect 31420 5940 31660 6180
rect 31750 5940 31990 6180
rect 32080 5940 32320 6180
rect 32410 5940 32650 6180
rect 32740 5940 32980 6180
rect 33070 5940 33310 6180
rect 33400 5940 33640 6180
rect 33730 5940 33970 6180
rect 34060 5940 34300 6180
rect 34390 5940 34630 6180
rect 34720 5940 34960 6180
rect 35050 5940 35290 6180
rect 28780 5610 29020 5850
rect 29110 5610 29350 5850
rect 29440 5610 29680 5850
rect 29770 5610 30010 5850
rect 30100 5610 30340 5850
rect 30430 5610 30670 5850
rect 30760 5610 31000 5850
rect 31090 5610 31330 5850
rect 31420 5610 31660 5850
rect 31750 5610 31990 5850
rect 32080 5610 32320 5850
rect 32410 5610 32650 5850
rect 32740 5610 32980 5850
rect 33070 5610 33310 5850
rect 33400 5610 33640 5850
rect 33730 5610 33970 5850
rect 34060 5610 34300 5850
rect 34390 5610 34630 5850
rect 34720 5610 34960 5850
rect 35050 5610 35290 5850
rect 28780 5280 29020 5520
rect 29110 5280 29350 5520
rect 29440 5280 29680 5520
rect 29770 5280 30010 5520
rect 30100 5280 30340 5520
rect 30430 5280 30670 5520
rect 30760 5280 31000 5520
rect 31090 5280 31330 5520
rect 31420 5280 31660 5520
rect 31750 5280 31990 5520
rect 32080 5280 32320 5520
rect 32410 5280 32650 5520
rect 32740 5280 32980 5520
rect 33070 5280 33310 5520
rect 33400 5280 33640 5520
rect 33730 5280 33970 5520
rect 34060 5280 34300 5520
rect 34390 5280 34630 5520
rect 34720 5280 34960 5520
rect 35050 5280 35290 5520
rect 28780 4950 29020 5190
rect 29110 4950 29350 5190
rect 29440 4950 29680 5190
rect 29770 4950 30010 5190
rect 30100 4950 30340 5190
rect 30430 4950 30670 5190
rect 30760 4950 31000 5190
rect 31090 4950 31330 5190
rect 31420 4950 31660 5190
rect 31750 4950 31990 5190
rect 32080 4950 32320 5190
rect 32410 4950 32650 5190
rect 32740 4950 32980 5190
rect 33070 4950 33310 5190
rect 33400 4950 33640 5190
rect 33730 4950 33970 5190
rect 34060 4950 34300 5190
rect 34390 4950 34630 5190
rect 34720 4950 34960 5190
rect 35050 4950 35290 5190
rect 28780 4620 29020 4860
rect 29110 4620 29350 4860
rect 29440 4620 29680 4860
rect 29770 4620 30010 4860
rect 30100 4620 30340 4860
rect 30430 4620 30670 4860
rect 30760 4620 31000 4860
rect 31090 4620 31330 4860
rect 31420 4620 31660 4860
rect 31750 4620 31990 4860
rect 32080 4620 32320 4860
rect 32410 4620 32650 4860
rect 32740 4620 32980 4860
rect 33070 4620 33310 4860
rect 33400 4620 33640 4860
rect 33730 4620 33970 4860
rect 34060 4620 34300 4860
rect 34390 4620 34630 4860
rect 34720 4620 34960 4860
rect 35050 4620 35290 4860
rect 28780 4290 29020 4530
rect 29110 4290 29350 4530
rect 29440 4290 29680 4530
rect 29770 4290 30010 4530
rect 30100 4290 30340 4530
rect 30430 4290 30670 4530
rect 30760 4290 31000 4530
rect 31090 4290 31330 4530
rect 31420 4290 31660 4530
rect 31750 4290 31990 4530
rect 32080 4290 32320 4530
rect 32410 4290 32650 4530
rect 32740 4290 32980 4530
rect 33070 4290 33310 4530
rect 33400 4290 33640 4530
rect 33730 4290 33970 4530
rect 34060 4290 34300 4530
rect 34390 4290 34630 4530
rect 34720 4290 34960 4530
rect 35050 4290 35290 4530
rect 28780 3960 29020 4200
rect 29110 3960 29350 4200
rect 29440 3960 29680 4200
rect 29770 3960 30010 4200
rect 30100 3960 30340 4200
rect 30430 3960 30670 4200
rect 30760 3960 31000 4200
rect 31090 3960 31330 4200
rect 31420 3960 31660 4200
rect 31750 3960 31990 4200
rect 32080 3960 32320 4200
rect 32410 3960 32650 4200
rect 32740 3960 32980 4200
rect 33070 3960 33310 4200
rect 33400 3960 33640 4200
rect 33730 3960 33970 4200
rect 34060 3960 34300 4200
rect 34390 3960 34630 4200
rect 34720 3960 34960 4200
rect 35050 3960 35290 4200
rect 28780 3630 29020 3870
rect 29110 3630 29350 3870
rect 29440 3630 29680 3870
rect 29770 3630 30010 3870
rect 30100 3630 30340 3870
rect 30430 3630 30670 3870
rect 30760 3630 31000 3870
rect 31090 3630 31330 3870
rect 31420 3630 31660 3870
rect 31750 3630 31990 3870
rect 32080 3630 32320 3870
rect 32410 3630 32650 3870
rect 32740 3630 32980 3870
rect 33070 3630 33310 3870
rect 33400 3630 33640 3870
rect 33730 3630 33970 3870
rect 34060 3630 34300 3870
rect 34390 3630 34630 3870
rect 34720 3630 34960 3870
rect 35050 3630 35290 3870
rect 28780 3300 29020 3540
rect 29110 3300 29350 3540
rect 29440 3300 29680 3540
rect 29770 3300 30010 3540
rect 30100 3300 30340 3540
rect 30430 3300 30670 3540
rect 30760 3300 31000 3540
rect 31090 3300 31330 3540
rect 31420 3300 31660 3540
rect 31750 3300 31990 3540
rect 32080 3300 32320 3540
rect 32410 3300 32650 3540
rect 32740 3300 32980 3540
rect 33070 3300 33310 3540
rect 33400 3300 33640 3540
rect 33730 3300 33970 3540
rect 34060 3300 34300 3540
rect 34390 3300 34630 3540
rect 34720 3300 34960 3540
rect 35050 3300 35290 3540
rect 28780 2970 29020 3210
rect 29110 2970 29350 3210
rect 29440 2970 29680 3210
rect 29770 2970 30010 3210
rect 30100 2970 30340 3210
rect 30430 2970 30670 3210
rect 30760 2970 31000 3210
rect 31090 2970 31330 3210
rect 31420 2970 31660 3210
rect 31750 2970 31990 3210
rect 32080 2970 32320 3210
rect 32410 2970 32650 3210
rect 32740 2970 32980 3210
rect 33070 2970 33310 3210
rect 33400 2970 33640 3210
rect 33730 2970 33970 3210
rect 34060 2970 34300 3210
rect 34390 2970 34630 3210
rect 34720 2970 34960 3210
rect 35050 2970 35290 3210
rect 28780 2640 29020 2880
rect 29110 2640 29350 2880
rect 29440 2640 29680 2880
rect 29770 2640 30010 2880
rect 30100 2640 30340 2880
rect 30430 2640 30670 2880
rect 30760 2640 31000 2880
rect 31090 2640 31330 2880
rect 31420 2640 31660 2880
rect 31750 2640 31990 2880
rect 32080 2640 32320 2880
rect 32410 2640 32650 2880
rect 32740 2640 32980 2880
rect 33070 2640 33310 2880
rect 33400 2640 33640 2880
rect 33730 2640 33970 2880
rect 34060 2640 34300 2880
rect 34390 2640 34630 2880
rect 34720 2640 34960 2880
rect 35050 2640 35290 2880
rect 28780 2310 29020 2550
rect 29110 2310 29350 2550
rect 29440 2310 29680 2550
rect 29770 2310 30010 2550
rect 30100 2310 30340 2550
rect 30430 2310 30670 2550
rect 30760 2310 31000 2550
rect 31090 2310 31330 2550
rect 31420 2310 31660 2550
rect 31750 2310 31990 2550
rect 32080 2310 32320 2550
rect 32410 2310 32650 2550
rect 32740 2310 32980 2550
rect 33070 2310 33310 2550
rect 33400 2310 33640 2550
rect 33730 2310 33970 2550
rect 34060 2310 34300 2550
rect 34390 2310 34630 2550
rect 34720 2310 34960 2550
rect 35050 2310 35290 2550
rect 28780 1980 29020 2220
rect 29110 1980 29350 2220
rect 29440 1980 29680 2220
rect 29770 1980 30010 2220
rect 30100 1980 30340 2220
rect 30430 1980 30670 2220
rect 30760 1980 31000 2220
rect 31090 1980 31330 2220
rect 31420 1980 31660 2220
rect 31750 1980 31990 2220
rect 32080 1980 32320 2220
rect 32410 1980 32650 2220
rect 32740 1980 32980 2220
rect 33070 1980 33310 2220
rect 33400 1980 33640 2220
rect 33730 1980 33970 2220
rect 34060 1980 34300 2220
rect 34390 1980 34630 2220
rect 34720 1980 34960 2220
rect 35050 1980 35290 2220
rect 28780 1650 29020 1890
rect 29110 1650 29350 1890
rect 29440 1650 29680 1890
rect 29770 1650 30010 1890
rect 30100 1650 30340 1890
rect 30430 1650 30670 1890
rect 30760 1650 31000 1890
rect 31090 1650 31330 1890
rect 31420 1650 31660 1890
rect 31750 1650 31990 1890
rect 32080 1650 32320 1890
rect 32410 1650 32650 1890
rect 32740 1650 32980 1890
rect 33070 1650 33310 1890
rect 33400 1650 33640 1890
rect 33730 1650 33970 1890
rect 34060 1650 34300 1890
rect 34390 1650 34630 1890
rect 34720 1650 34960 1890
rect 35050 1650 35290 1890
rect 28780 1320 29020 1560
rect 29110 1320 29350 1560
rect 29440 1320 29680 1560
rect 29770 1320 30010 1560
rect 30100 1320 30340 1560
rect 30430 1320 30670 1560
rect 30760 1320 31000 1560
rect 31090 1320 31330 1560
rect 31420 1320 31660 1560
rect 31750 1320 31990 1560
rect 32080 1320 32320 1560
rect 32410 1320 32650 1560
rect 32740 1320 32980 1560
rect 33070 1320 33310 1560
rect 33400 1320 33640 1560
rect 33730 1320 33970 1560
rect 34060 1320 34300 1560
rect 34390 1320 34630 1560
rect 34720 1320 34960 1560
rect 35050 1320 35290 1560
rect 28780 -10 29020 230
rect 29110 -10 29350 230
rect 29440 -10 29680 230
rect 29770 -10 30010 230
rect 30100 -10 30340 230
rect 30430 -10 30670 230
rect 30760 -10 31000 230
rect 31090 -10 31330 230
rect 31420 -10 31660 230
rect 31750 -10 31990 230
rect 32080 -10 32320 230
rect 32410 -10 32650 230
rect 32740 -10 32980 230
rect 33070 -10 33310 230
rect 33400 -10 33640 230
rect 33730 -10 33970 230
rect 34060 -10 34300 230
rect 34390 -10 34630 230
rect 34720 -10 34960 230
rect 35050 -10 35290 230
rect 28780 -340 29020 -100
rect 29110 -340 29350 -100
rect 29440 -340 29680 -100
rect 29770 -340 30010 -100
rect 30100 -340 30340 -100
rect 30430 -340 30670 -100
rect 30760 -340 31000 -100
rect 31090 -340 31330 -100
rect 31420 -340 31660 -100
rect 31750 -340 31990 -100
rect 32080 -340 32320 -100
rect 32410 -340 32650 -100
rect 32740 -340 32980 -100
rect 33070 -340 33310 -100
rect 33400 -340 33640 -100
rect 33730 -340 33970 -100
rect 34060 -340 34300 -100
rect 34390 -340 34630 -100
rect 34720 -340 34960 -100
rect 35050 -340 35290 -100
rect 28780 -670 29020 -430
rect 29110 -670 29350 -430
rect 29440 -670 29680 -430
rect 29770 -670 30010 -430
rect 30100 -670 30340 -430
rect 30430 -670 30670 -430
rect 30760 -670 31000 -430
rect 31090 -670 31330 -430
rect 31420 -670 31660 -430
rect 31750 -670 31990 -430
rect 32080 -670 32320 -430
rect 32410 -670 32650 -430
rect 32740 -670 32980 -430
rect 33070 -670 33310 -430
rect 33400 -670 33640 -430
rect 33730 -670 33970 -430
rect 34060 -670 34300 -430
rect 34390 -670 34630 -430
rect 34720 -670 34960 -430
rect 35050 -670 35290 -430
rect 28780 -1000 29020 -760
rect 29110 -1000 29350 -760
rect 29440 -1000 29680 -760
rect 29770 -1000 30010 -760
rect 30100 -1000 30340 -760
rect 30430 -1000 30670 -760
rect 30760 -1000 31000 -760
rect 31090 -1000 31330 -760
rect 31420 -1000 31660 -760
rect 31750 -1000 31990 -760
rect 32080 -1000 32320 -760
rect 32410 -1000 32650 -760
rect 32740 -1000 32980 -760
rect 33070 -1000 33310 -760
rect 33400 -1000 33640 -760
rect 33730 -1000 33970 -760
rect 34060 -1000 34300 -760
rect 34390 -1000 34630 -760
rect 34720 -1000 34960 -760
rect 35050 -1000 35290 -760
rect 28780 -1330 29020 -1090
rect 29110 -1330 29350 -1090
rect 29440 -1330 29680 -1090
rect 29770 -1330 30010 -1090
rect 30100 -1330 30340 -1090
rect 30430 -1330 30670 -1090
rect 30760 -1330 31000 -1090
rect 31090 -1330 31330 -1090
rect 31420 -1330 31660 -1090
rect 31750 -1330 31990 -1090
rect 32080 -1330 32320 -1090
rect 32410 -1330 32650 -1090
rect 32740 -1330 32980 -1090
rect 33070 -1330 33310 -1090
rect 33400 -1330 33640 -1090
rect 33730 -1330 33970 -1090
rect 34060 -1330 34300 -1090
rect 34390 -1330 34630 -1090
rect 34720 -1330 34960 -1090
rect 35050 -1330 35290 -1090
rect 28780 -1660 29020 -1420
rect 29110 -1660 29350 -1420
rect 29440 -1660 29680 -1420
rect 29770 -1660 30010 -1420
rect 30100 -1660 30340 -1420
rect 30430 -1660 30670 -1420
rect 30760 -1660 31000 -1420
rect 31090 -1660 31330 -1420
rect 31420 -1660 31660 -1420
rect 31750 -1660 31990 -1420
rect 32080 -1660 32320 -1420
rect 32410 -1660 32650 -1420
rect 32740 -1660 32980 -1420
rect 33070 -1660 33310 -1420
rect 33400 -1660 33640 -1420
rect 33730 -1660 33970 -1420
rect 34060 -1660 34300 -1420
rect 34390 -1660 34630 -1420
rect 34720 -1660 34960 -1420
rect 35050 -1660 35290 -1420
rect 28780 -1990 29020 -1750
rect 29110 -1990 29350 -1750
rect 29440 -1990 29680 -1750
rect 29770 -1990 30010 -1750
rect 30100 -1990 30340 -1750
rect 30430 -1990 30670 -1750
rect 30760 -1990 31000 -1750
rect 31090 -1990 31330 -1750
rect 31420 -1990 31660 -1750
rect 31750 -1990 31990 -1750
rect 32080 -1990 32320 -1750
rect 32410 -1990 32650 -1750
rect 32740 -1990 32980 -1750
rect 33070 -1990 33310 -1750
rect 33400 -1990 33640 -1750
rect 33730 -1990 33970 -1750
rect 34060 -1990 34300 -1750
rect 34390 -1990 34630 -1750
rect 34720 -1990 34960 -1750
rect 35050 -1990 35290 -1750
rect 28780 -2320 29020 -2080
rect 29110 -2320 29350 -2080
rect 29440 -2320 29680 -2080
rect 29770 -2320 30010 -2080
rect 30100 -2320 30340 -2080
rect 30430 -2320 30670 -2080
rect 30760 -2320 31000 -2080
rect 31090 -2320 31330 -2080
rect 31420 -2320 31660 -2080
rect 31750 -2320 31990 -2080
rect 32080 -2320 32320 -2080
rect 32410 -2320 32650 -2080
rect 32740 -2320 32980 -2080
rect 33070 -2320 33310 -2080
rect 33400 -2320 33640 -2080
rect 33730 -2320 33970 -2080
rect 34060 -2320 34300 -2080
rect 34390 -2320 34630 -2080
rect 34720 -2320 34960 -2080
rect 35050 -2320 35290 -2080
rect 28780 -2650 29020 -2410
rect 29110 -2650 29350 -2410
rect 29440 -2650 29680 -2410
rect 29770 -2650 30010 -2410
rect 30100 -2650 30340 -2410
rect 30430 -2650 30670 -2410
rect 30760 -2650 31000 -2410
rect 31090 -2650 31330 -2410
rect 31420 -2650 31660 -2410
rect 31750 -2650 31990 -2410
rect 32080 -2650 32320 -2410
rect 32410 -2650 32650 -2410
rect 32740 -2650 32980 -2410
rect 33070 -2650 33310 -2410
rect 33400 -2650 33640 -2410
rect 33730 -2650 33970 -2410
rect 34060 -2650 34300 -2410
rect 34390 -2650 34630 -2410
rect 34720 -2650 34960 -2410
rect 35050 -2650 35290 -2410
rect 28780 -2980 29020 -2740
rect 29110 -2980 29350 -2740
rect 29440 -2980 29680 -2740
rect 29770 -2980 30010 -2740
rect 30100 -2980 30340 -2740
rect 30430 -2980 30670 -2740
rect 30760 -2980 31000 -2740
rect 31090 -2980 31330 -2740
rect 31420 -2980 31660 -2740
rect 31750 -2980 31990 -2740
rect 32080 -2980 32320 -2740
rect 32410 -2980 32650 -2740
rect 32740 -2980 32980 -2740
rect 33070 -2980 33310 -2740
rect 33400 -2980 33640 -2740
rect 33730 -2980 33970 -2740
rect 34060 -2980 34300 -2740
rect 34390 -2980 34630 -2740
rect 34720 -2980 34960 -2740
rect 35050 -2980 35290 -2740
rect 28780 -3310 29020 -3070
rect 29110 -3310 29350 -3070
rect 29440 -3310 29680 -3070
rect 29770 -3310 30010 -3070
rect 30100 -3310 30340 -3070
rect 30430 -3310 30670 -3070
rect 30760 -3310 31000 -3070
rect 31090 -3310 31330 -3070
rect 31420 -3310 31660 -3070
rect 31750 -3310 31990 -3070
rect 32080 -3310 32320 -3070
rect 32410 -3310 32650 -3070
rect 32740 -3310 32980 -3070
rect 33070 -3310 33310 -3070
rect 33400 -3310 33640 -3070
rect 33730 -3310 33970 -3070
rect 34060 -3310 34300 -3070
rect 34390 -3310 34630 -3070
rect 34720 -3310 34960 -3070
rect 35050 -3310 35290 -3070
rect 28780 -3640 29020 -3400
rect 29110 -3640 29350 -3400
rect 29440 -3640 29680 -3400
rect 29770 -3640 30010 -3400
rect 30100 -3640 30340 -3400
rect 30430 -3640 30670 -3400
rect 30760 -3640 31000 -3400
rect 31090 -3640 31330 -3400
rect 31420 -3640 31660 -3400
rect 31750 -3640 31990 -3400
rect 32080 -3640 32320 -3400
rect 32410 -3640 32650 -3400
rect 32740 -3640 32980 -3400
rect 33070 -3640 33310 -3400
rect 33400 -3640 33640 -3400
rect 33730 -3640 33970 -3400
rect 34060 -3640 34300 -3400
rect 34390 -3640 34630 -3400
rect 34720 -3640 34960 -3400
rect 35050 -3640 35290 -3400
rect 28780 -3970 29020 -3730
rect 29110 -3970 29350 -3730
rect 29440 -3970 29680 -3730
rect 29770 -3970 30010 -3730
rect 30100 -3970 30340 -3730
rect 30430 -3970 30670 -3730
rect 30760 -3970 31000 -3730
rect 31090 -3970 31330 -3730
rect 31420 -3970 31660 -3730
rect 31750 -3970 31990 -3730
rect 32080 -3970 32320 -3730
rect 32410 -3970 32650 -3730
rect 32740 -3970 32980 -3730
rect 33070 -3970 33310 -3730
rect 33400 -3970 33640 -3730
rect 33730 -3970 33970 -3730
rect 34060 -3970 34300 -3730
rect 34390 -3970 34630 -3730
rect 34720 -3970 34960 -3730
rect 35050 -3970 35290 -3730
rect -1650 -4500 -1410 -4260
rect -1320 -4500 -1080 -4260
rect -990 -4500 -750 -4260
rect -660 -4500 -420 -4260
rect -1650 -4830 -1410 -4590
rect -1320 -4830 -1080 -4590
rect -990 -4830 -750 -4590
rect -660 -4830 -420 -4590
rect -1650 -5160 -1410 -4920
rect -1320 -5160 -1080 -4920
rect -990 -5160 -750 -4920
rect -660 -5160 -420 -4920
rect -1650 -5490 -1410 -5250
rect -1320 -5490 -1080 -5250
rect -990 -5490 -750 -5250
rect -660 -5490 -420 -5250
rect 28780 -4300 29020 -4060
rect 29110 -4300 29350 -4060
rect 29440 -4300 29680 -4060
rect 29770 -4300 30010 -4060
rect 30100 -4300 30340 -4060
rect 30430 -4300 30670 -4060
rect 30760 -4300 31000 -4060
rect 31090 -4300 31330 -4060
rect 31420 -4300 31660 -4060
rect 31750 -4300 31990 -4060
rect 32080 -4300 32320 -4060
rect 32410 -4300 32650 -4060
rect 32740 -4300 32980 -4060
rect 33070 -4300 33310 -4060
rect 33400 -4300 33640 -4060
rect 33730 -4300 33970 -4060
rect 34060 -4300 34300 -4060
rect 34390 -4300 34630 -4060
rect 34720 -4300 34960 -4060
rect 35050 -4300 35290 -4060
rect 28780 -4630 29020 -4390
rect 29110 -4630 29350 -4390
rect 29440 -4630 29680 -4390
rect 29770 -4630 30010 -4390
rect 30100 -4630 30340 -4390
rect 30430 -4630 30670 -4390
rect 30760 -4630 31000 -4390
rect 31090 -4630 31330 -4390
rect 31420 -4630 31660 -4390
rect 31750 -4630 31990 -4390
rect 32080 -4630 32320 -4390
rect 32410 -4630 32650 -4390
rect 32740 -4630 32980 -4390
rect 33070 -4630 33310 -4390
rect 33400 -4630 33640 -4390
rect 33730 -4630 33970 -4390
rect 34060 -4630 34300 -4390
rect 34390 -4630 34630 -4390
rect 34720 -4630 34960 -4390
rect 35050 -4630 35290 -4390
rect 28780 -4960 29020 -4720
rect 29110 -4960 29350 -4720
rect 29440 -4960 29680 -4720
rect 29770 -4960 30010 -4720
rect 30100 -4960 30340 -4720
rect 30430 -4960 30670 -4720
rect 30760 -4960 31000 -4720
rect 31090 -4960 31330 -4720
rect 31420 -4960 31660 -4720
rect 31750 -4960 31990 -4720
rect 32080 -4960 32320 -4720
rect 32410 -4960 32650 -4720
rect 32740 -4960 32980 -4720
rect 33070 -4960 33310 -4720
rect 33400 -4960 33640 -4720
rect 33730 -4960 33970 -4720
rect 34060 -4960 34300 -4720
rect 34390 -4960 34630 -4720
rect 34720 -4960 34960 -4720
rect 35050 -4960 35290 -4720
rect 28780 -5290 29020 -5050
rect 29110 -5290 29350 -5050
rect 29440 -5290 29680 -5050
rect 29770 -5290 30010 -5050
rect 30100 -5290 30340 -5050
rect 30430 -5290 30670 -5050
rect 30760 -5290 31000 -5050
rect 31090 -5290 31330 -5050
rect 31420 -5290 31660 -5050
rect 31750 -5290 31990 -5050
rect 32080 -5290 32320 -5050
rect 32410 -5290 32650 -5050
rect 32740 -5290 32980 -5050
rect 33070 -5290 33310 -5050
rect 33400 -5290 33640 -5050
rect 33730 -5290 33970 -5050
rect 34060 -5290 34300 -5050
rect 34390 -5290 34630 -5050
rect 34720 -5290 34960 -5050
rect 35050 -5290 35290 -5050
rect 28780 -5620 29020 -5380
rect 29110 -5620 29350 -5380
rect 29440 -5620 29680 -5380
rect 29770 -5620 30010 -5380
rect 30100 -5620 30340 -5380
rect 30430 -5620 30670 -5380
rect 30760 -5620 31000 -5380
rect 31090 -5620 31330 -5380
rect 31420 -5620 31660 -5380
rect 31750 -5620 31990 -5380
rect 32080 -5620 32320 -5380
rect 32410 -5620 32650 -5380
rect 32740 -5620 32980 -5380
rect 33070 -5620 33310 -5380
rect 33400 -5620 33640 -5380
rect 33730 -5620 33970 -5380
rect 34060 -5620 34300 -5380
rect 34390 -5620 34630 -5380
rect 34720 -5620 34960 -5380
rect 35050 -5620 35290 -5380
rect 28780 -5950 29020 -5710
rect 29110 -5950 29350 -5710
rect 29440 -5950 29680 -5710
rect 29770 -5950 30010 -5710
rect 30100 -5950 30340 -5710
rect 30430 -5950 30670 -5710
rect 30760 -5950 31000 -5710
rect 31090 -5950 31330 -5710
rect 31420 -5950 31660 -5710
rect 31750 -5950 31990 -5710
rect 32080 -5950 32320 -5710
rect 32410 -5950 32650 -5710
rect 32740 -5950 32980 -5710
rect 33070 -5950 33310 -5710
rect 33400 -5950 33640 -5710
rect 33730 -5950 33970 -5710
rect 34060 -5950 34300 -5710
rect 34390 -5950 34630 -5710
rect 34720 -5950 34960 -5710
rect 35050 -5950 35290 -5710
rect 28780 -6280 29020 -6040
rect 29110 -6280 29350 -6040
rect 29440 -6280 29680 -6040
rect 29770 -6280 30010 -6040
rect 30100 -6280 30340 -6040
rect 30430 -6280 30670 -6040
rect 30760 -6280 31000 -6040
rect 31090 -6280 31330 -6040
rect 31420 -6280 31660 -6040
rect 31750 -6280 31990 -6040
rect 32080 -6280 32320 -6040
rect 32410 -6280 32650 -6040
rect 32740 -6280 32980 -6040
rect 33070 -6280 33310 -6040
rect 33400 -6280 33640 -6040
rect 33730 -6280 33970 -6040
rect 34060 -6280 34300 -6040
rect 34390 -6280 34630 -6040
rect 34720 -6280 34960 -6040
rect 35050 -6280 35290 -6040
rect -1650 -7900 -1410 -7660
rect -1320 -7900 -1080 -7660
rect -990 -7900 -750 -7660
rect -660 -7900 -420 -7660
rect -1650 -8230 -1410 -7990
rect -1320 -8230 -1080 -7990
rect -990 -8230 -750 -7990
rect -660 -8230 -420 -7990
rect -1650 -8560 -1410 -8320
rect -1320 -8560 -1080 -8320
rect -990 -8560 -750 -8320
rect -660 -8560 -420 -8320
rect -1650 -8890 -1410 -8650
rect -1320 -8890 -1080 -8650
rect -990 -8890 -750 -8650
rect -660 -8890 -420 -8650
<< metal5 >>
rect -5020 20790 7290 21140
rect -5020 20550 -4670 20790
rect -4430 20550 -4340 20790
rect -4100 20550 -4010 20790
rect -3770 20550 -3680 20790
rect -3440 20550 -3350 20790
rect -3110 20550 -3020 20790
rect -2780 20550 -2690 20790
rect -2450 20550 -2360 20790
rect -2120 20550 -2030 20790
rect -1790 20550 -1700 20790
rect -1460 20550 -1370 20790
rect -1130 20550 -1040 20790
rect -800 20550 -710 20790
rect -470 20550 -380 20790
rect -140 20550 -50 20790
rect 190 20550 280 20790
rect 520 20550 610 20790
rect 850 20550 940 20790
rect 1180 20550 1270 20790
rect 1510 20550 1600 20790
rect 1840 20550 1930 20790
rect 2170 20550 2260 20790
rect 2500 20550 2590 20790
rect 2830 20550 2920 20790
rect 3160 20550 3250 20790
rect 3490 20550 3580 20790
rect 3820 20550 3910 20790
rect 4150 20550 4240 20790
rect 4480 20550 4570 20790
rect 4810 20550 4900 20790
rect 5140 20550 5230 20790
rect 5470 20550 5560 20790
rect 5800 20550 5890 20790
rect 6130 20550 6220 20790
rect 6460 20550 6550 20790
rect 6790 20550 6880 20790
rect 7120 20550 7290 20790
rect -5020 20460 7290 20550
rect -5020 20220 -4670 20460
rect -4430 20220 -4340 20460
rect -4100 20220 -4010 20460
rect -3770 20220 -3680 20460
rect -3440 20220 -3350 20460
rect -3110 20220 -3020 20460
rect -2780 20220 -2690 20460
rect -2450 20220 -2360 20460
rect -2120 20220 -2030 20460
rect -1790 20220 -1700 20460
rect -1460 20220 -1370 20460
rect -1130 20220 -1040 20460
rect -800 20220 -710 20460
rect -470 20220 -380 20460
rect -140 20220 -50 20460
rect 190 20220 280 20460
rect 520 20220 610 20460
rect 850 20220 940 20460
rect 1180 20220 1270 20460
rect 1510 20220 1600 20460
rect 1840 20220 1930 20460
rect 2170 20220 2260 20460
rect 2500 20220 2590 20460
rect 2830 20220 2920 20460
rect 3160 20220 3250 20460
rect 3490 20220 3580 20460
rect 3820 20220 3910 20460
rect 4150 20220 4240 20460
rect 4480 20220 4570 20460
rect 4810 20220 4900 20460
rect 5140 20220 5230 20460
rect 5470 20220 5560 20460
rect 5800 20220 5890 20460
rect 6130 20220 6220 20460
rect 6460 20220 6550 20460
rect 6790 20220 6880 20460
rect 7120 20220 7290 20460
rect -5020 20130 7290 20220
rect -5020 19890 -4670 20130
rect -4430 19890 -4340 20130
rect -4100 19890 -4010 20130
rect -3770 19890 -3680 20130
rect -3440 19890 -3350 20130
rect -3110 19890 -3020 20130
rect -2780 19890 -2690 20130
rect -2450 19890 -2360 20130
rect -2120 19890 -2030 20130
rect -1790 19890 -1700 20130
rect -1460 19890 -1370 20130
rect -1130 19890 -1040 20130
rect -800 19890 -710 20130
rect -470 19890 -380 20130
rect -140 19890 -50 20130
rect 190 19890 280 20130
rect 520 19890 610 20130
rect 850 19890 940 20130
rect 1180 19890 1270 20130
rect 1510 19890 1600 20130
rect 1840 19890 1930 20130
rect 2170 19890 2260 20130
rect 2500 19890 2590 20130
rect 2830 19890 2920 20130
rect 3160 19890 3250 20130
rect 3490 19890 3580 20130
rect 3820 19890 3910 20130
rect 4150 19890 4240 20130
rect 4480 19890 4570 20130
rect 4810 19890 4900 20130
rect 5140 19890 5230 20130
rect 5470 19890 5560 20130
rect 5800 19890 5890 20130
rect 6130 19890 6220 20130
rect 6460 19890 6550 20130
rect 6790 19890 6880 20130
rect 7120 19890 7290 20130
rect -5020 19800 7290 19890
rect -5020 19560 -4670 19800
rect -4430 19560 -4340 19800
rect -4100 19560 -4010 19800
rect -3770 19560 -3680 19800
rect -3440 19560 -3350 19800
rect -3110 19560 -3020 19800
rect -2780 19560 -2690 19800
rect -2450 19560 -2360 19800
rect -2120 19560 -2030 19800
rect -1790 19560 -1700 19800
rect -1460 19560 -1370 19800
rect -1130 19560 -1040 19800
rect -800 19560 -710 19800
rect -470 19560 -380 19800
rect -140 19560 -50 19800
rect 190 19560 280 19800
rect 520 19560 610 19800
rect 850 19560 940 19800
rect 1180 19560 1270 19800
rect 1510 19560 1600 19800
rect 1840 19560 1930 19800
rect 2170 19560 2260 19800
rect 2500 19560 2590 19800
rect 2830 19560 2920 19800
rect 3160 19560 3250 19800
rect 3490 19560 3580 19800
rect 3820 19560 3910 19800
rect 4150 19560 4240 19800
rect 4480 19560 4570 19800
rect 4810 19560 4900 19800
rect 5140 19560 5230 19800
rect 5470 19560 5560 19800
rect 5800 19560 5890 19800
rect 6130 19560 6220 19800
rect 6460 19560 6550 19800
rect 6790 19560 6880 19800
rect 7120 19560 7290 19800
rect -5020 19470 7290 19560
rect -5020 19230 -4670 19470
rect -4430 19230 -4340 19470
rect -4100 19230 -4010 19470
rect -3770 19230 -3680 19470
rect -3440 19230 -3350 19470
rect -3110 19230 -3020 19470
rect -2780 19230 -2690 19470
rect -2450 19230 -2360 19470
rect -2120 19230 -2030 19470
rect -1790 19230 -1700 19470
rect -1460 19230 -1370 19470
rect -1130 19230 -1040 19470
rect -800 19230 -710 19470
rect -470 19230 -380 19470
rect -140 19230 -50 19470
rect 190 19230 280 19470
rect 520 19230 610 19470
rect 850 19230 940 19470
rect 1180 19230 1270 19470
rect 1510 19230 1600 19470
rect 1840 19230 1930 19470
rect 2170 19230 2260 19470
rect 2500 19230 2590 19470
rect 2830 19230 2920 19470
rect 3160 19230 3250 19470
rect 3490 19230 3580 19470
rect 3820 19230 3910 19470
rect 4150 19230 4240 19470
rect 4480 19230 4570 19470
rect 4810 19230 4900 19470
rect 5140 19230 5230 19470
rect 5470 19230 5560 19470
rect 5800 19230 5890 19470
rect 6130 19230 6220 19470
rect 6460 19230 6550 19470
rect 6790 19230 6880 19470
rect 7120 19230 7290 19470
rect -5020 19140 7290 19230
rect -5020 18900 -4670 19140
rect -4430 18900 -4340 19140
rect -4100 18900 -4010 19140
rect -3770 18900 -3680 19140
rect -3440 18900 -3350 19140
rect -3110 18900 -3020 19140
rect -2780 18900 -2690 19140
rect -2450 18900 -2360 19140
rect -2120 18900 -2030 19140
rect -1790 18900 -1700 19140
rect -1460 18900 -1370 19140
rect -1130 18900 -1040 19140
rect -800 18900 -710 19140
rect -470 18900 -380 19140
rect -140 18900 -50 19140
rect 190 18900 280 19140
rect 520 18900 610 19140
rect 850 18900 940 19140
rect 1180 18900 1270 19140
rect 1510 18900 1600 19140
rect 1840 18900 1930 19140
rect 2170 18900 2260 19140
rect 2500 18900 2590 19140
rect 2830 18900 2920 19140
rect 3160 18900 3250 19140
rect 3490 18900 3580 19140
rect 3820 18900 3910 19140
rect 4150 18900 4240 19140
rect 4480 18900 4570 19140
rect 4810 18900 4900 19140
rect 5140 18900 5230 19140
rect 5470 18900 5560 19140
rect 5800 18900 5890 19140
rect 6130 18900 6220 19140
rect 6460 18900 6550 19140
rect 6790 18900 6880 19140
rect 7120 18900 7290 19140
rect -5020 18810 7290 18900
rect -5020 18570 -4670 18810
rect -4430 18570 -4340 18810
rect -4100 18570 -4010 18810
rect -3770 18570 -3680 18810
rect -3440 18570 -3350 18810
rect -3110 18570 -3020 18810
rect -2780 18570 -2690 18810
rect -2450 18570 -2360 18810
rect -2120 18570 -2030 18810
rect -1790 18570 -1700 18810
rect -1460 18570 -1370 18810
rect -1130 18570 -1040 18810
rect -800 18570 -710 18810
rect -470 18570 -380 18810
rect -140 18570 -50 18810
rect 190 18570 280 18810
rect 520 18570 610 18810
rect 850 18570 940 18810
rect 1180 18570 1270 18810
rect 1510 18570 1600 18810
rect 1840 18570 1930 18810
rect 2170 18570 2260 18810
rect 2500 18570 2590 18810
rect 2830 18570 2920 18810
rect 3160 18570 3250 18810
rect 3490 18570 3580 18810
rect 3820 18570 3910 18810
rect 4150 18570 4240 18810
rect 4480 18570 4570 18810
rect 4810 18570 4900 18810
rect 5140 18570 5230 18810
rect 5470 18570 5560 18810
rect 5800 18570 5890 18810
rect 6130 18570 6220 18810
rect 6460 18570 6550 18810
rect 6790 18570 6880 18810
rect 7120 18570 7290 18810
rect -5020 18480 7290 18570
rect -5020 18240 -4670 18480
rect -4430 18240 -4340 18480
rect -4100 18240 -4010 18480
rect -3770 18240 -3680 18480
rect -3440 18240 -3350 18480
rect -3110 18240 -3020 18480
rect -2780 18240 -2690 18480
rect -2450 18240 -2360 18480
rect -2120 18240 -2030 18480
rect -1790 18240 -1700 18480
rect -1460 18240 -1370 18480
rect -1130 18240 -1040 18480
rect -800 18240 -710 18480
rect -470 18240 -380 18480
rect -140 18240 -50 18480
rect 190 18240 280 18480
rect 520 18240 610 18480
rect 850 18240 940 18480
rect 1180 18240 1270 18480
rect 1510 18240 1600 18480
rect 1840 18240 1930 18480
rect 2170 18240 2260 18480
rect 2500 18240 2590 18480
rect 2830 18240 2920 18480
rect 3160 18240 3250 18480
rect 3490 18240 3580 18480
rect 3820 18240 3910 18480
rect 4150 18240 4240 18480
rect 4480 18240 4570 18480
rect 4810 18240 4900 18480
rect 5140 18240 5230 18480
rect 5470 18240 5560 18480
rect 5800 18240 5890 18480
rect 6130 18240 6220 18480
rect 6460 18240 6550 18480
rect 6790 18240 6880 18480
rect 7120 18240 7290 18480
rect -5020 18150 7290 18240
rect -5020 17910 -4670 18150
rect -4430 17910 -4340 18150
rect -4100 17910 -4010 18150
rect -3770 17910 -3680 18150
rect -3440 17910 -3350 18150
rect -3110 17910 -3020 18150
rect -2780 17910 -2690 18150
rect -2450 17910 -2360 18150
rect -2120 17910 -2030 18150
rect -1790 17910 -1700 18150
rect -1460 17910 -1370 18150
rect -1130 17910 -1040 18150
rect -800 17910 -710 18150
rect -470 17910 -380 18150
rect -140 17910 -50 18150
rect 190 17910 280 18150
rect 520 17910 610 18150
rect 850 17910 940 18150
rect 1180 17910 1270 18150
rect 1510 17910 1600 18150
rect 1840 17910 1930 18150
rect 2170 17910 2260 18150
rect 2500 17910 2590 18150
rect 2830 17910 2920 18150
rect 3160 17910 3250 18150
rect 3490 17910 3580 18150
rect 3820 17910 3910 18150
rect 4150 17910 4240 18150
rect 4480 17910 4570 18150
rect 4810 17910 4900 18150
rect 5140 17910 5230 18150
rect 5470 17910 5560 18150
rect 5800 17910 5890 18150
rect 6130 17910 6220 18150
rect 6460 17910 6550 18150
rect 6790 17910 6880 18150
rect 7120 17910 7290 18150
rect -5020 17820 7290 17910
rect -5020 17580 -4670 17820
rect -4430 17580 -4340 17820
rect -4100 17580 -4010 17820
rect -3770 17580 -3680 17820
rect -3440 17580 -3350 17820
rect -3110 17580 -3020 17820
rect -2780 17580 -2690 17820
rect -2450 17580 -2360 17820
rect -2120 17580 -2030 17820
rect -1790 17580 -1700 17820
rect -1460 17580 -1370 17820
rect -1130 17580 -1040 17820
rect -800 17580 -710 17820
rect -470 17580 -380 17820
rect -140 17580 -50 17820
rect 190 17580 280 17820
rect 520 17580 610 17820
rect 850 17580 940 17820
rect 1180 17580 1270 17820
rect 1510 17580 1600 17820
rect 1840 17580 1930 17820
rect 2170 17580 2260 17820
rect 2500 17580 2590 17820
rect 2830 17580 2920 17820
rect 3160 17580 3250 17820
rect 3490 17580 3580 17820
rect 3820 17580 3910 17820
rect 4150 17580 4240 17820
rect 4480 17580 4570 17820
rect 4810 17580 4900 17820
rect 5140 17580 5230 17820
rect 5470 17580 5560 17820
rect 5800 17580 5890 17820
rect 6130 17580 6220 17820
rect 6460 17580 6550 17820
rect 6790 17580 6880 17820
rect 7120 17580 7290 17820
rect -5020 17490 7290 17580
rect -5020 17250 -4670 17490
rect -4430 17250 -4340 17490
rect -4100 17250 -4010 17490
rect -3770 17250 -3680 17490
rect -3440 17250 -3350 17490
rect -3110 17250 -3020 17490
rect -2780 17250 -2690 17490
rect -2450 17250 -2360 17490
rect -2120 17250 -2030 17490
rect -1790 17250 -1700 17490
rect -1460 17250 -1370 17490
rect -1130 17250 -1040 17490
rect -800 17250 -710 17490
rect -470 17250 -380 17490
rect -140 17250 -50 17490
rect 190 17250 280 17490
rect 520 17250 610 17490
rect 850 17250 940 17490
rect 1180 17250 1270 17490
rect 1510 17250 1600 17490
rect 1840 17250 1930 17490
rect 2170 17250 2260 17490
rect 2500 17250 2590 17490
rect 2830 17250 2920 17490
rect 3160 17250 3250 17490
rect 3490 17250 3580 17490
rect 3820 17250 3910 17490
rect 4150 17250 4240 17490
rect 4480 17250 4570 17490
rect 4810 17250 4900 17490
rect 5140 17250 5230 17490
rect 5470 17250 5560 17490
rect 5800 17250 5890 17490
rect 6130 17250 6220 17490
rect 6460 17250 6550 17490
rect 6790 17250 6880 17490
rect 7120 17250 7290 17490
rect -5020 17160 7290 17250
rect -5020 16920 -4670 17160
rect -4430 16920 -4340 17160
rect -4100 16920 -4010 17160
rect -3770 16920 -3680 17160
rect -3440 16920 -3350 17160
rect -3110 16920 -3020 17160
rect -2780 16920 -2690 17160
rect -2450 16920 -2360 17160
rect -2120 16920 -2030 17160
rect -1790 16920 -1700 17160
rect -1460 16920 -1370 17160
rect -1130 16920 -1040 17160
rect -800 16920 -710 17160
rect -470 16920 -380 17160
rect -140 16920 -50 17160
rect 190 16920 280 17160
rect 520 16920 610 17160
rect 850 16920 940 17160
rect 1180 16920 1270 17160
rect 1510 16920 1600 17160
rect 1840 16920 1930 17160
rect 2170 16920 2260 17160
rect 2500 16920 2590 17160
rect 2830 16920 2920 17160
rect 3160 16920 3250 17160
rect 3490 16920 3580 17160
rect 3820 16920 3910 17160
rect 4150 16920 4240 17160
rect 4480 16920 4570 17160
rect 4810 16920 4900 17160
rect 5140 16920 5230 17160
rect 5470 16920 5560 17160
rect 5800 16920 5890 17160
rect 6130 16920 6220 17160
rect 6460 16920 6550 17160
rect 6790 16920 6880 17160
rect 7120 16920 7290 17160
rect -5020 16830 7290 16920
rect -5020 16590 -4670 16830
rect -4430 16590 -4340 16830
rect -4100 16590 -4010 16830
rect -3770 16590 -3680 16830
rect -3440 16590 -3350 16830
rect -3110 16590 -3020 16830
rect -2780 16590 -2690 16830
rect -2450 16590 -2360 16830
rect -2120 16590 -2030 16830
rect -1790 16590 -1700 16830
rect -1460 16590 -1370 16830
rect -1130 16590 -1040 16830
rect -800 16590 -710 16830
rect -470 16590 -380 16830
rect -140 16590 -50 16830
rect 190 16590 280 16830
rect 520 16590 610 16830
rect 850 16590 940 16830
rect 1180 16590 1270 16830
rect 1510 16590 1600 16830
rect 1840 16590 1930 16830
rect 2170 16590 2260 16830
rect 2500 16590 2590 16830
rect 2830 16590 2920 16830
rect 3160 16590 3250 16830
rect 3490 16590 3580 16830
rect 3820 16590 3910 16830
rect 4150 16590 4240 16830
rect 4480 16590 4570 16830
rect 4810 16590 4900 16830
rect 5140 16590 5230 16830
rect 5470 16590 5560 16830
rect 5800 16590 5890 16830
rect 6130 16590 6220 16830
rect 6460 16590 6550 16830
rect 6790 16590 6880 16830
rect 7120 16590 7290 16830
rect -5020 16500 7290 16590
rect -5020 16260 -4670 16500
rect -4430 16260 -4340 16500
rect -4100 16260 -4010 16500
rect -3770 16260 -3680 16500
rect -3440 16260 -3350 16500
rect -3110 16260 -3020 16500
rect -2780 16260 -2690 16500
rect -2450 16260 -2360 16500
rect -2120 16260 -2030 16500
rect -1790 16260 -1700 16500
rect -1460 16260 -1370 16500
rect -1130 16260 -1040 16500
rect -800 16260 -710 16500
rect -470 16260 -380 16500
rect -140 16260 -50 16500
rect 190 16260 280 16500
rect 520 16260 610 16500
rect 850 16260 940 16500
rect 1180 16260 1270 16500
rect 1510 16260 1600 16500
rect 1840 16260 1930 16500
rect 2170 16260 2260 16500
rect 2500 16260 2590 16500
rect 2830 16260 2920 16500
rect 3160 16260 3250 16500
rect 3490 16260 3580 16500
rect 3820 16260 3910 16500
rect 4150 16260 4240 16500
rect 4480 16260 4570 16500
rect 4810 16260 4900 16500
rect 5140 16260 5230 16500
rect 5470 16260 5560 16500
rect 5800 16260 5890 16500
rect 6130 16260 6220 16500
rect 6460 16260 6550 16500
rect 6790 16260 6880 16500
rect 7120 16260 7290 16500
rect -5020 16170 7290 16260
rect -5020 15930 -4670 16170
rect -4430 15930 -4340 16170
rect -4100 15930 -4010 16170
rect -3770 15930 -3680 16170
rect -3440 15930 -3350 16170
rect -3110 15930 -3020 16170
rect -2780 15930 -2690 16170
rect -2450 15930 -2360 16170
rect -2120 15930 -2030 16170
rect -1790 15930 -1700 16170
rect -1460 15930 -1370 16170
rect -1130 15930 -1040 16170
rect -800 15930 -710 16170
rect -470 15930 -380 16170
rect -140 15930 -50 16170
rect 190 15930 280 16170
rect 520 15930 610 16170
rect 850 15930 940 16170
rect 1180 15930 1270 16170
rect 1510 15930 1600 16170
rect 1840 15930 1930 16170
rect 2170 15930 2260 16170
rect 2500 15930 2590 16170
rect 2830 15930 2920 16170
rect 3160 15930 3250 16170
rect 3490 15930 3580 16170
rect 3820 15930 3910 16170
rect 4150 15930 4240 16170
rect 4480 15930 4570 16170
rect 4810 15930 4900 16170
rect 5140 15930 5230 16170
rect 5470 15930 5560 16170
rect 5800 15930 5890 16170
rect 6130 15930 6220 16170
rect 6460 15930 6550 16170
rect 6790 15930 6880 16170
rect 7120 15930 7290 16170
rect -5020 15840 7290 15930
rect -5020 15600 -4670 15840
rect -4430 15600 -4340 15840
rect -4100 15600 -4010 15840
rect -3770 15600 -3680 15840
rect -3440 15600 -3350 15840
rect -3110 15600 -3020 15840
rect -2780 15600 -2690 15840
rect -2450 15600 -2360 15840
rect -2120 15600 -2030 15840
rect -1790 15600 -1700 15840
rect -1460 15600 -1370 15840
rect -1130 15600 -1040 15840
rect -800 15600 -710 15840
rect -470 15600 -380 15840
rect -140 15600 -50 15840
rect 190 15600 280 15840
rect 520 15600 610 15840
rect 850 15600 940 15840
rect 1180 15600 1270 15840
rect 1510 15600 1600 15840
rect 1840 15600 1930 15840
rect 2170 15600 2260 15840
rect 2500 15600 2590 15840
rect 2830 15600 2920 15840
rect 3160 15600 3250 15840
rect 3490 15600 3580 15840
rect 3820 15600 3910 15840
rect 4150 15600 4240 15840
rect 4480 15600 4570 15840
rect 4810 15600 4900 15840
rect 5140 15600 5230 15840
rect 5470 15600 5560 15840
rect 5800 15600 5890 15840
rect 6130 15600 6220 15840
rect 6460 15600 6550 15840
rect 6790 15600 6880 15840
rect 7120 15600 7290 15840
rect -5020 15510 7290 15600
rect -5020 15270 -4670 15510
rect -4430 15270 -4340 15510
rect -4100 15270 -4010 15510
rect -3770 15270 -3680 15510
rect -3440 15270 -3350 15510
rect -3110 15270 -3020 15510
rect -2780 15270 -2690 15510
rect -2450 15270 -2360 15510
rect -2120 15270 -2030 15510
rect -1790 15270 -1700 15510
rect -1460 15270 -1370 15510
rect -1130 15270 -1040 15510
rect -800 15270 -710 15510
rect -470 15270 -380 15510
rect -140 15270 -50 15510
rect 190 15270 280 15510
rect 520 15270 610 15510
rect 850 15270 940 15510
rect 1180 15270 1270 15510
rect 1510 15270 1600 15510
rect 1840 15270 1930 15510
rect 2170 15270 2260 15510
rect 2500 15270 2590 15510
rect 2830 15270 2920 15510
rect 3160 15270 3250 15510
rect 3490 15270 3580 15510
rect 3820 15270 3910 15510
rect 4150 15270 4240 15510
rect 4480 15270 4570 15510
rect 4810 15270 4900 15510
rect 5140 15270 5230 15510
rect 5470 15270 5560 15510
rect 5800 15270 5890 15510
rect 6130 15270 6220 15510
rect 6460 15270 6550 15510
rect 6790 15270 6880 15510
rect 7120 15270 7290 15510
rect -5020 15180 7290 15270
rect -5020 14940 -4670 15180
rect -4430 14940 -4340 15180
rect -4100 14940 -4010 15180
rect -3770 14940 -3680 15180
rect -3440 14940 -3350 15180
rect -3110 14940 -3020 15180
rect -2780 14940 -2690 15180
rect -2450 14940 -2360 15180
rect -2120 14940 -2030 15180
rect -1790 14940 -1700 15180
rect -1460 14940 -1370 15180
rect -1130 14940 -1040 15180
rect -800 14940 -710 15180
rect -470 14940 -380 15180
rect -140 14940 -50 15180
rect 190 14940 280 15180
rect 520 14940 610 15180
rect 850 14940 940 15180
rect 1180 14940 1270 15180
rect 1510 14940 1600 15180
rect 1840 14940 1930 15180
rect 2170 14940 2260 15180
rect 2500 14940 2590 15180
rect 2830 14940 2920 15180
rect 3160 14940 3250 15180
rect 3490 14940 3580 15180
rect 3820 14940 3910 15180
rect 4150 14940 4240 15180
rect 4480 14940 4570 15180
rect 4810 14940 4900 15180
rect 5140 14940 5230 15180
rect 5470 14940 5560 15180
rect 5800 14940 5890 15180
rect 6130 14940 6220 15180
rect 6460 14940 6550 15180
rect 6790 14940 6880 15180
rect 7120 14940 7290 15180
rect -5020 14850 7290 14940
rect -5020 14610 -4670 14850
rect -4430 14610 -4340 14850
rect -4100 14610 -4010 14850
rect -3770 14610 -3680 14850
rect -3440 14610 -3350 14850
rect -3110 14610 -3020 14850
rect -2780 14610 -2690 14850
rect -2450 14610 -2360 14850
rect -2120 14610 -2030 14850
rect -1790 14610 -1700 14850
rect -1460 14610 -1370 14850
rect -1130 14610 -1040 14850
rect -800 14610 -710 14850
rect -470 14610 -380 14850
rect -140 14610 -50 14850
rect 190 14610 280 14850
rect 520 14610 610 14850
rect 850 14610 940 14850
rect 1180 14610 1270 14850
rect 1510 14610 1600 14850
rect 1840 14610 1930 14850
rect 2170 14610 2260 14850
rect 2500 14610 2590 14850
rect 2830 14610 2920 14850
rect 3160 14610 3250 14850
rect 3490 14610 3580 14850
rect 3820 14610 3910 14850
rect 4150 14610 4240 14850
rect 4480 14610 4570 14850
rect 4810 14610 4900 14850
rect 5140 14610 5230 14850
rect 5470 14610 5560 14850
rect 5800 14610 5890 14850
rect 6130 14610 6220 14850
rect 6460 14610 6550 14850
rect 6790 14610 6880 14850
rect 7120 14610 7290 14850
rect -5020 14520 7290 14610
rect -5020 14280 -4670 14520
rect -4430 14280 -4340 14520
rect -4100 14280 -4010 14520
rect -3770 14280 -3680 14520
rect -3440 14280 -3350 14520
rect -3110 14280 -3020 14520
rect -2780 14280 -2690 14520
rect -2450 14280 -2360 14520
rect -2120 14280 -2030 14520
rect -1790 14280 -1700 14520
rect -1460 14280 -1370 14520
rect -1130 14280 -1040 14520
rect -800 14280 -710 14520
rect -470 14280 -380 14520
rect -140 14280 -50 14520
rect 190 14280 280 14520
rect 520 14280 610 14520
rect 850 14280 940 14520
rect 1180 14280 1270 14520
rect 1510 14280 1600 14520
rect 1840 14280 1930 14520
rect 2170 14280 2260 14520
rect 2500 14280 2590 14520
rect 2830 14280 2920 14520
rect 3160 14280 3250 14520
rect 3490 14280 3580 14520
rect 3820 14280 3910 14520
rect 4150 14280 4240 14520
rect 4480 14280 4570 14520
rect 4810 14280 4900 14520
rect 5140 14280 5230 14520
rect 5470 14280 5560 14520
rect 5800 14280 5890 14520
rect 6130 14280 6220 14520
rect 6460 14280 6550 14520
rect 6790 14280 6880 14520
rect 7120 14280 7290 14520
rect -5020 14190 7290 14280
rect -5020 13950 -4670 14190
rect -4430 13950 -4340 14190
rect -4100 13950 -4010 14190
rect -3770 13950 -3680 14190
rect -3440 13950 -3350 14190
rect -3110 13950 -3020 14190
rect -2780 13950 -2690 14190
rect -2450 13950 -2360 14190
rect -2120 13950 -2030 14190
rect -1790 13950 -1700 14190
rect -1460 13950 -1370 14190
rect -1130 13950 -1040 14190
rect -800 13950 -710 14190
rect -470 13950 -380 14190
rect -140 13950 -50 14190
rect 190 13950 280 14190
rect 520 13950 610 14190
rect 850 13950 940 14190
rect 1180 13950 1270 14190
rect 1510 13950 1600 14190
rect 1840 13950 1930 14190
rect 2170 13950 2260 14190
rect 2500 13950 2590 14190
rect 2830 13950 2920 14190
rect 3160 13950 3250 14190
rect 3490 13950 3580 14190
rect 3820 13950 3910 14190
rect 4150 13950 4240 14190
rect 4480 13950 4570 14190
rect 4810 13950 4900 14190
rect 5140 13950 5230 14190
rect 5470 13950 5560 14190
rect 5800 13950 5890 14190
rect 6130 13950 6220 14190
rect 6460 13950 6550 14190
rect 6790 13950 6880 14190
rect 7120 13950 7290 14190
rect -5020 13860 7290 13950
rect -5020 13620 -4670 13860
rect -4430 13620 -4340 13860
rect -4100 13620 -4010 13860
rect -3770 13620 -3680 13860
rect -3440 13620 -3350 13860
rect -3110 13620 -3020 13860
rect -2780 13620 -2690 13860
rect -2450 13620 -2360 13860
rect -2120 13620 -2030 13860
rect -1790 13620 -1700 13860
rect -1460 13620 -1370 13860
rect -1130 13620 -1040 13860
rect -800 13620 -710 13860
rect -470 13620 -380 13860
rect -140 13620 -50 13860
rect 190 13620 280 13860
rect 520 13620 610 13860
rect 850 13620 940 13860
rect 1180 13620 1270 13860
rect 1510 13620 1600 13860
rect 1840 13620 1930 13860
rect 2170 13620 2260 13860
rect 2500 13620 2590 13860
rect 2830 13620 2920 13860
rect 3160 13620 3250 13860
rect 3490 13620 3580 13860
rect 3820 13620 3910 13860
rect 4150 13620 4240 13860
rect 4480 13620 4570 13860
rect 4810 13620 4900 13860
rect 5140 13620 5230 13860
rect 5470 13620 5560 13860
rect 5800 13620 5890 13860
rect 6130 13620 6220 13860
rect 6460 13620 6550 13860
rect 6790 13620 6880 13860
rect 7120 13620 7290 13860
rect -5020 13530 7290 13620
rect -5020 13290 -4670 13530
rect -4430 13290 -4340 13530
rect -4100 13290 -4010 13530
rect -3770 13290 -3680 13530
rect -3440 13290 -3350 13530
rect -3110 13290 -3020 13530
rect -2780 13290 -2690 13530
rect -2450 13290 -2360 13530
rect -2120 13290 -2030 13530
rect -1790 13290 -1700 13530
rect -1460 13290 -1370 13530
rect -1130 13290 -1040 13530
rect -800 13290 -710 13530
rect -470 13290 -380 13530
rect -140 13290 -50 13530
rect 190 13290 280 13530
rect 520 13290 610 13530
rect 850 13290 940 13530
rect 1180 13290 1270 13530
rect 1510 13290 1600 13530
rect 1840 13290 1930 13530
rect 2170 13290 2260 13530
rect 2500 13290 2590 13530
rect 2830 13290 2920 13530
rect 3160 13290 3250 13530
rect 3490 13290 3580 13530
rect 3820 13290 3910 13530
rect 4150 13290 4240 13530
rect 4480 13290 4570 13530
rect 4810 13290 4900 13530
rect 5140 13290 5230 13530
rect 5470 13290 5560 13530
rect 5800 13290 5890 13530
rect 6130 13290 6220 13530
rect 6460 13290 6550 13530
rect 6790 13290 6880 13530
rect 7120 13290 7290 13530
rect -5020 13200 7290 13290
rect -5020 12960 -4670 13200
rect -4430 12960 -4340 13200
rect -4100 12960 -4010 13200
rect -3770 12960 -3680 13200
rect -3440 12960 -3350 13200
rect -3110 12960 -3020 13200
rect -2780 12960 -2690 13200
rect -2450 12960 -2360 13200
rect -2120 12960 -2030 13200
rect -1790 12960 -1700 13200
rect -1460 12960 -1370 13200
rect -1130 12960 -1040 13200
rect -800 12960 -710 13200
rect -470 12960 -380 13200
rect -140 12960 -50 13200
rect 190 12960 280 13200
rect 520 12960 610 13200
rect 850 12960 940 13200
rect 1180 12960 1270 13200
rect 1510 12960 1600 13200
rect 1840 12960 1930 13200
rect 2170 12960 2260 13200
rect 2500 12960 2590 13200
rect 2830 12960 2920 13200
rect 3160 12960 3250 13200
rect 3490 12960 3580 13200
rect 3820 12960 3910 13200
rect 4150 12960 4240 13200
rect 4480 12960 4570 13200
rect 4810 12960 4900 13200
rect 5140 12960 5230 13200
rect 5470 12960 5560 13200
rect 5800 12960 5890 13200
rect 6130 12960 6220 13200
rect 6460 12960 6550 13200
rect 6790 12960 6880 13200
rect 7120 12960 7290 13200
rect -5020 12870 7290 12960
rect -5020 12630 -4670 12870
rect -4430 12630 -4340 12870
rect -4100 12630 -4010 12870
rect -3770 12630 -3680 12870
rect -3440 12630 -3350 12870
rect -3110 12630 -3020 12870
rect -2780 12630 -2690 12870
rect -2450 12630 -2360 12870
rect -2120 12630 -2030 12870
rect -1790 12630 -1700 12870
rect -1460 12630 -1370 12870
rect -1130 12630 -1040 12870
rect -800 12630 -710 12870
rect -470 12630 -380 12870
rect -140 12630 -50 12870
rect 190 12630 280 12870
rect 520 12630 610 12870
rect 850 12630 940 12870
rect 1180 12630 1270 12870
rect 1510 12630 1600 12870
rect 1840 12630 1930 12870
rect 2170 12630 2260 12870
rect 2500 12630 2590 12870
rect 2830 12630 2920 12870
rect 3160 12630 3250 12870
rect 3490 12630 3580 12870
rect 3820 12630 3910 12870
rect 4150 12630 4240 12870
rect 4480 12630 4570 12870
rect 4810 12630 4900 12870
rect 5140 12630 5230 12870
rect 5470 12630 5560 12870
rect 5800 12630 5890 12870
rect 6130 12630 6220 12870
rect 6460 12630 6550 12870
rect 6790 12630 6880 12870
rect 7120 12630 7290 12870
rect -5020 12540 7290 12630
rect -5020 12300 -4670 12540
rect -4430 12300 -4340 12540
rect -4100 12300 -4010 12540
rect -3770 12300 -3680 12540
rect -3440 12300 -3350 12540
rect -3110 12300 -3020 12540
rect -2780 12300 -2690 12540
rect -2450 12300 -2360 12540
rect -2120 12300 -2030 12540
rect -1790 12300 -1700 12540
rect -1460 12300 -1370 12540
rect -1130 12300 -1040 12540
rect -800 12300 -710 12540
rect -470 12300 -380 12540
rect -140 12300 -50 12540
rect 190 12300 280 12540
rect 520 12300 610 12540
rect 850 12300 940 12540
rect 1180 12300 1270 12540
rect 1510 12300 1600 12540
rect 1840 12300 1930 12540
rect 2170 12300 2260 12540
rect 2500 12300 2590 12540
rect 2830 12300 2920 12540
rect 3160 12300 3250 12540
rect 3490 12300 3580 12540
rect 3820 12300 3910 12540
rect 4150 12300 4240 12540
rect 4480 12300 4570 12540
rect 4810 12300 4900 12540
rect 5140 12300 5230 12540
rect 5470 12300 5560 12540
rect 5800 12300 5890 12540
rect 6130 12300 6220 12540
rect 6460 12300 6550 12540
rect 6790 12300 6880 12540
rect 7120 12300 7290 12540
rect -5020 12210 7290 12300
rect -5020 11970 -4670 12210
rect -4430 11970 -4340 12210
rect -4100 11970 -4010 12210
rect -3770 11970 -3680 12210
rect -3440 11970 -3350 12210
rect -3110 11970 -3020 12210
rect -2780 11970 -2690 12210
rect -2450 11970 -2360 12210
rect -2120 11970 -2030 12210
rect -1790 11970 -1700 12210
rect -1460 11970 -1370 12210
rect -1130 11970 -1040 12210
rect -800 11970 -710 12210
rect -470 11970 -380 12210
rect -140 11970 -50 12210
rect 190 11970 280 12210
rect 520 11970 610 12210
rect 850 11970 940 12210
rect 1180 11970 1270 12210
rect 1510 11970 1600 12210
rect 1840 11970 1930 12210
rect 2170 11970 2260 12210
rect 2500 11970 2590 12210
rect 2830 11970 2920 12210
rect 3160 11970 3250 12210
rect 3490 11970 3580 12210
rect 3820 11970 3910 12210
rect 4150 11970 4240 12210
rect 4480 11970 4570 12210
rect 4810 11970 4900 12210
rect 5140 11970 5230 12210
rect 5470 11970 5560 12210
rect 5800 11970 5890 12210
rect 6130 11970 6220 12210
rect 6460 11970 6550 12210
rect 6790 11970 6880 12210
rect 7120 11970 7290 12210
rect -5020 11880 7290 11970
rect -5020 11640 -4670 11880
rect -4430 11640 -4340 11880
rect -4100 11640 -4010 11880
rect -3770 11640 -3680 11880
rect -3440 11640 -3350 11880
rect -3110 11640 -3020 11880
rect -2780 11640 -2690 11880
rect -2450 11640 -2360 11880
rect -2120 11640 -2030 11880
rect -1790 11640 -1700 11880
rect -1460 11640 -1370 11880
rect -1130 11640 -1040 11880
rect -800 11640 -710 11880
rect -470 11640 -380 11880
rect -140 11640 -50 11880
rect 190 11640 280 11880
rect 520 11640 610 11880
rect 850 11640 940 11880
rect 1180 11640 1270 11880
rect 1510 11640 1600 11880
rect 1840 11640 1930 11880
rect 2170 11640 2260 11880
rect 2500 11640 2590 11880
rect 2830 11640 2920 11880
rect 3160 11640 3250 11880
rect 3490 11640 3580 11880
rect 3820 11640 3910 11880
rect 4150 11640 4240 11880
rect 4480 11640 4570 11880
rect 4810 11640 4900 11880
rect 5140 11640 5230 11880
rect 5470 11640 5560 11880
rect 5800 11640 5890 11880
rect 6130 11640 6220 11880
rect 6460 11640 6550 11880
rect 6790 11640 6880 11880
rect 7120 11640 7290 11880
rect -5020 11550 7290 11640
rect -5020 11310 -4670 11550
rect -4430 11310 -4340 11550
rect -4100 11310 -4010 11550
rect -3770 11310 -3680 11550
rect -3440 11310 -3350 11550
rect -3110 11310 -3020 11550
rect -2780 11310 -2690 11550
rect -2450 11310 -2360 11550
rect -2120 11310 -2030 11550
rect -1790 11310 -1700 11550
rect -1460 11310 -1370 11550
rect -1130 11310 -1040 11550
rect -800 11310 -710 11550
rect -470 11310 -380 11550
rect -140 11310 -50 11550
rect 190 11310 280 11550
rect 520 11310 610 11550
rect 850 11310 940 11550
rect 1180 11310 1270 11550
rect 1510 11310 1600 11550
rect 1840 11310 1930 11550
rect 2170 11310 2260 11550
rect 2500 11310 2590 11550
rect 2830 11310 2920 11550
rect 3160 11310 3250 11550
rect 3490 11310 3580 11550
rect 3820 11310 3910 11550
rect 4150 11310 4240 11550
rect 4480 11310 4570 11550
rect 4810 11310 4900 11550
rect 5140 11310 5230 11550
rect 5470 11310 5560 11550
rect 5800 11310 5890 11550
rect 6130 11310 6220 11550
rect 6460 11310 6550 11550
rect 6790 11310 6880 11550
rect 7120 11310 7290 11550
rect -5020 11220 7290 11310
rect -5020 10980 -4670 11220
rect -4430 10980 -4340 11220
rect -4100 10980 -4010 11220
rect -3770 10980 -3680 11220
rect -3440 10980 -3350 11220
rect -3110 10980 -3020 11220
rect -2780 10980 -2690 11220
rect -2450 10980 -2360 11220
rect -2120 10980 -2030 11220
rect -1790 10980 -1700 11220
rect -1460 10980 -1370 11220
rect -1130 10980 -1040 11220
rect -800 10980 -710 11220
rect -470 10980 -380 11220
rect -140 10980 -50 11220
rect 190 10980 280 11220
rect 520 10980 610 11220
rect 850 10980 940 11220
rect 1180 10980 1270 11220
rect 1510 10980 1600 11220
rect 1840 10980 1930 11220
rect 2170 10980 2260 11220
rect 2500 10980 2590 11220
rect 2830 10980 2920 11220
rect 3160 10980 3250 11220
rect 3490 10980 3580 11220
rect 3820 10980 3910 11220
rect 4150 10980 4240 11220
rect 4480 10980 4570 11220
rect 4810 10980 4900 11220
rect 5140 10980 5230 11220
rect 5470 10980 5560 11220
rect 5800 10980 5890 11220
rect 6130 10980 6220 11220
rect 6460 10980 6550 11220
rect 6790 10980 6880 11220
rect 7120 10980 7290 11220
rect -5020 10890 7290 10980
rect -5020 10650 -4670 10890
rect -4430 10650 -4340 10890
rect -4100 10650 -4010 10890
rect -3770 10650 -3680 10890
rect -3440 10650 -3350 10890
rect -3110 10650 -3020 10890
rect -2780 10650 -2690 10890
rect -2450 10650 -2360 10890
rect -2120 10650 -2030 10890
rect -1790 10650 -1700 10890
rect -1460 10650 -1370 10890
rect -1130 10650 -1040 10890
rect -800 10650 -710 10890
rect -470 10650 -380 10890
rect -140 10650 -50 10890
rect 190 10650 280 10890
rect 520 10650 610 10890
rect 850 10650 940 10890
rect 1180 10650 1270 10890
rect 1510 10650 1600 10890
rect 1840 10650 1930 10890
rect 2170 10650 2260 10890
rect 2500 10650 2590 10890
rect 2830 10650 2920 10890
rect 3160 10650 3250 10890
rect 3490 10650 3580 10890
rect 3820 10650 3910 10890
rect 4150 10650 4240 10890
rect 4480 10650 4570 10890
rect 4810 10650 4900 10890
rect 5140 10650 5230 10890
rect 5470 10650 5560 10890
rect 5800 10650 5890 10890
rect 6130 10650 6220 10890
rect 6460 10650 6550 10890
rect 6790 10650 6880 10890
rect 7120 10650 7290 10890
rect -5020 10560 7290 10650
rect -5020 10320 -4670 10560
rect -4430 10320 -4340 10560
rect -4100 10320 -4010 10560
rect -3770 10320 -3680 10560
rect -3440 10320 -3350 10560
rect -3110 10320 -3020 10560
rect -2780 10320 -2690 10560
rect -2450 10320 -2360 10560
rect -2120 10320 -2030 10560
rect -1790 10320 -1700 10560
rect -1460 10320 -1370 10560
rect -1130 10320 -1040 10560
rect -800 10320 -710 10560
rect -470 10320 -380 10560
rect -140 10320 -50 10560
rect 190 10320 280 10560
rect 520 10320 610 10560
rect 850 10320 940 10560
rect 1180 10320 1270 10560
rect 1510 10320 1600 10560
rect 1840 10320 1930 10560
rect 2170 10320 2260 10560
rect 2500 10320 2590 10560
rect 2830 10320 2920 10560
rect 3160 10320 3250 10560
rect 3490 10320 3580 10560
rect 3820 10320 3910 10560
rect 4150 10320 4240 10560
rect 4480 10320 4570 10560
rect 4810 10320 4900 10560
rect 5140 10320 5230 10560
rect 5470 10320 5560 10560
rect 5800 10320 5890 10560
rect 6130 10320 6220 10560
rect 6460 10320 6550 10560
rect 6790 10320 6880 10560
rect 7120 10320 7290 10560
rect -5020 10230 7290 10320
rect -5020 9990 -4670 10230
rect -4430 9990 -4340 10230
rect -4100 9990 -4010 10230
rect -3770 9990 -3680 10230
rect -3440 9990 -3350 10230
rect -3110 9990 -3020 10230
rect -2780 9990 -2690 10230
rect -2450 9990 -2360 10230
rect -2120 9990 -2030 10230
rect -1790 9990 -1700 10230
rect -1460 9990 -1370 10230
rect -1130 9990 -1040 10230
rect -800 9990 -710 10230
rect -470 9990 -380 10230
rect -140 9990 -50 10230
rect 190 9990 280 10230
rect 520 9990 610 10230
rect 850 9990 940 10230
rect 1180 9990 1270 10230
rect 1510 9990 1600 10230
rect 1840 9990 1930 10230
rect 2170 9990 2260 10230
rect 2500 9990 2590 10230
rect 2830 9990 2920 10230
rect 3160 9990 3250 10230
rect 3490 9990 3580 10230
rect 3820 9990 3910 10230
rect 4150 9990 4240 10230
rect 4480 9990 4570 10230
rect 4810 9990 4900 10230
rect 5140 9990 5230 10230
rect 5470 9990 5560 10230
rect 5800 9990 5890 10230
rect 6130 9990 6220 10230
rect 6460 9990 6550 10230
rect 6790 9990 6880 10230
rect 7120 9990 7290 10230
rect -5020 9900 7290 9990
rect -5020 9660 -4670 9900
rect -4430 9660 -4340 9900
rect -4100 9660 -4010 9900
rect -3770 9660 -3680 9900
rect -3440 9660 -3350 9900
rect -3110 9660 -3020 9900
rect -2780 9660 -2690 9900
rect -2450 9660 -2360 9900
rect -2120 9660 -2030 9900
rect -1790 9660 -1700 9900
rect -1460 9660 -1370 9900
rect -1130 9660 -1040 9900
rect -800 9660 -710 9900
rect -470 9660 -380 9900
rect -140 9660 -50 9900
rect 190 9660 280 9900
rect 520 9660 610 9900
rect 850 9660 940 9900
rect 1180 9660 1270 9900
rect 1510 9660 1600 9900
rect 1840 9660 1930 9900
rect 2170 9660 2260 9900
rect 2500 9660 2590 9900
rect 2830 9660 2920 9900
rect 3160 9660 3250 9900
rect 3490 9660 3580 9900
rect 3820 9660 3910 9900
rect 4150 9660 4240 9900
rect 4480 9660 4570 9900
rect 4810 9660 4900 9900
rect 5140 9660 5230 9900
rect 5470 9660 5560 9900
rect 5800 9660 5890 9900
rect 6130 9660 6220 9900
rect 6460 9660 6550 9900
rect 6790 9660 6880 9900
rect 7120 9660 7290 9900
rect -5020 9570 7290 9660
rect -5020 9330 -4670 9570
rect -4430 9330 -4340 9570
rect -4100 9330 -4010 9570
rect -3770 9330 -3680 9570
rect -3440 9330 -3350 9570
rect -3110 9330 -3020 9570
rect -2780 9330 -2690 9570
rect -2450 9330 -2360 9570
rect -2120 9330 -2030 9570
rect -1790 9330 -1700 9570
rect -1460 9330 -1370 9570
rect -1130 9330 -1040 9570
rect -800 9330 -710 9570
rect -470 9330 -380 9570
rect -140 9330 -50 9570
rect 190 9330 280 9570
rect 520 9330 610 9570
rect 850 9330 940 9570
rect 1180 9330 1270 9570
rect 1510 9330 1600 9570
rect 1840 9330 1930 9570
rect 2170 9330 2260 9570
rect 2500 9330 2590 9570
rect 2830 9330 2920 9570
rect 3160 9330 3250 9570
rect 3490 9330 3580 9570
rect 3820 9330 3910 9570
rect 4150 9330 4240 9570
rect 4480 9330 4570 9570
rect 4810 9330 4900 9570
rect 5140 9330 5230 9570
rect 5470 9330 5560 9570
rect 5800 9330 5890 9570
rect 6130 9330 6220 9570
rect 6460 9330 6550 9570
rect 6790 9330 6880 9570
rect 7120 9330 7290 9570
rect -5020 9240 7290 9330
rect -5020 9000 -4670 9240
rect -4430 9000 -4340 9240
rect -4100 9000 -4010 9240
rect -3770 9000 -3680 9240
rect -3440 9000 -3350 9240
rect -3110 9000 -3020 9240
rect -2780 9000 -2690 9240
rect -2450 9000 -2360 9240
rect -2120 9000 -2030 9240
rect -1790 9000 -1700 9240
rect -1460 9000 -1370 9240
rect -1130 9000 -1040 9240
rect -800 9000 -710 9240
rect -470 9000 -380 9240
rect -140 9000 -50 9240
rect 190 9000 280 9240
rect 520 9000 610 9240
rect 850 9000 940 9240
rect 1180 9000 1270 9240
rect 1510 9000 1600 9240
rect 1840 9000 1930 9240
rect 2170 9000 2260 9240
rect 2500 9000 2590 9240
rect 2830 9000 2920 9240
rect 3160 9000 3250 9240
rect 3490 9000 3580 9240
rect 3820 9000 3910 9240
rect 4150 9000 4240 9240
rect 4480 9000 4570 9240
rect 4810 9000 4900 9240
rect 5140 9000 5230 9240
rect 5470 9000 5560 9240
rect 5800 9000 5890 9240
rect 6130 9000 6220 9240
rect 6460 9000 6550 9240
rect 6790 9000 6880 9240
rect 7120 9000 7290 9240
rect -5020 8460 7290 9000
rect -5020 8220 -4650 8460
rect -4410 8220 -4320 8460
rect -4080 8220 -3990 8460
rect -3750 8220 -3660 8460
rect -3420 8220 -3330 8460
rect -3090 8220 -3000 8460
rect -2760 8220 -2670 8460
rect -2430 8220 -2340 8460
rect -2100 8220 -2010 8460
rect -1770 8220 -1640 8460
rect -1400 8220 -1310 8460
rect -1070 8220 -980 8460
rect -740 8220 -650 8460
rect -410 8220 -320 8460
rect -80 8220 10 8460
rect 250 8220 340 8460
rect 580 8220 670 8460
rect 910 8220 1000 8460
rect 1240 8220 1370 8460
rect 1610 8220 1700 8460
rect 1940 8220 2030 8460
rect 2270 8220 2360 8460
rect 2600 8220 2690 8460
rect 2930 8220 3020 8460
rect 3260 8220 3350 8460
rect 3590 8220 3680 8460
rect 3920 8220 4010 8460
rect 4250 8220 4380 8460
rect 4620 8220 4710 8460
rect 4950 8220 5040 8460
rect 5280 8220 5370 8460
rect 5610 8220 5700 8460
rect 5940 8220 6030 8460
rect 6270 8220 6360 8460
rect 6600 8220 6690 8460
rect 6930 8220 7020 8460
rect 7260 8220 7290 8460
rect -5020 8190 7290 8220
rect 7610 20790 19920 21140
rect 7610 20550 7780 20790
rect 8020 20550 8110 20790
rect 8350 20550 8440 20790
rect 8680 20550 8770 20790
rect 9010 20550 9100 20790
rect 9340 20550 9430 20790
rect 9670 20550 9760 20790
rect 10000 20550 10090 20790
rect 10330 20550 10420 20790
rect 10660 20550 10750 20790
rect 10990 20550 11080 20790
rect 11320 20550 11410 20790
rect 11650 20550 11740 20790
rect 11980 20550 12070 20790
rect 12310 20550 12400 20790
rect 12640 20550 12730 20790
rect 12970 20550 13060 20790
rect 13300 20550 13390 20790
rect 13630 20550 13720 20790
rect 13960 20550 14050 20790
rect 14290 20550 14380 20790
rect 14620 20550 14710 20790
rect 14950 20550 15040 20790
rect 15280 20550 15370 20790
rect 15610 20550 15700 20790
rect 15940 20550 16030 20790
rect 16270 20550 16360 20790
rect 16600 20550 16690 20790
rect 16930 20550 17020 20790
rect 17260 20550 17350 20790
rect 17590 20550 17680 20790
rect 17920 20550 18010 20790
rect 18250 20550 18340 20790
rect 18580 20550 18670 20790
rect 18910 20550 19000 20790
rect 19240 20550 19330 20790
rect 19570 20550 19920 20790
rect 7610 20460 19920 20550
rect 7610 20220 7780 20460
rect 8020 20220 8110 20460
rect 8350 20220 8440 20460
rect 8680 20220 8770 20460
rect 9010 20220 9100 20460
rect 9340 20220 9430 20460
rect 9670 20220 9760 20460
rect 10000 20220 10090 20460
rect 10330 20220 10420 20460
rect 10660 20220 10750 20460
rect 10990 20220 11080 20460
rect 11320 20220 11410 20460
rect 11650 20220 11740 20460
rect 11980 20220 12070 20460
rect 12310 20220 12400 20460
rect 12640 20220 12730 20460
rect 12970 20220 13060 20460
rect 13300 20220 13390 20460
rect 13630 20220 13720 20460
rect 13960 20220 14050 20460
rect 14290 20220 14380 20460
rect 14620 20220 14710 20460
rect 14950 20220 15040 20460
rect 15280 20220 15370 20460
rect 15610 20220 15700 20460
rect 15940 20220 16030 20460
rect 16270 20220 16360 20460
rect 16600 20220 16690 20460
rect 16930 20220 17020 20460
rect 17260 20220 17350 20460
rect 17590 20220 17680 20460
rect 17920 20220 18010 20460
rect 18250 20220 18340 20460
rect 18580 20220 18670 20460
rect 18910 20220 19000 20460
rect 19240 20220 19330 20460
rect 19570 20220 19920 20460
rect 7610 20130 19920 20220
rect 7610 19890 7780 20130
rect 8020 19890 8110 20130
rect 8350 19890 8440 20130
rect 8680 19890 8770 20130
rect 9010 19890 9100 20130
rect 9340 19890 9430 20130
rect 9670 19890 9760 20130
rect 10000 19890 10090 20130
rect 10330 19890 10420 20130
rect 10660 19890 10750 20130
rect 10990 19890 11080 20130
rect 11320 19890 11410 20130
rect 11650 19890 11740 20130
rect 11980 19890 12070 20130
rect 12310 19890 12400 20130
rect 12640 19890 12730 20130
rect 12970 19890 13060 20130
rect 13300 19890 13390 20130
rect 13630 19890 13720 20130
rect 13960 19890 14050 20130
rect 14290 19890 14380 20130
rect 14620 19890 14710 20130
rect 14950 19890 15040 20130
rect 15280 19890 15370 20130
rect 15610 19890 15700 20130
rect 15940 19890 16030 20130
rect 16270 19890 16360 20130
rect 16600 19890 16690 20130
rect 16930 19890 17020 20130
rect 17260 19890 17350 20130
rect 17590 19890 17680 20130
rect 17920 19890 18010 20130
rect 18250 19890 18340 20130
rect 18580 19890 18670 20130
rect 18910 19890 19000 20130
rect 19240 19890 19330 20130
rect 19570 19890 19920 20130
rect 7610 19800 19920 19890
rect 7610 19560 7780 19800
rect 8020 19560 8110 19800
rect 8350 19560 8440 19800
rect 8680 19560 8770 19800
rect 9010 19560 9100 19800
rect 9340 19560 9430 19800
rect 9670 19560 9760 19800
rect 10000 19560 10090 19800
rect 10330 19560 10420 19800
rect 10660 19560 10750 19800
rect 10990 19560 11080 19800
rect 11320 19560 11410 19800
rect 11650 19560 11740 19800
rect 11980 19560 12070 19800
rect 12310 19560 12400 19800
rect 12640 19560 12730 19800
rect 12970 19560 13060 19800
rect 13300 19560 13390 19800
rect 13630 19560 13720 19800
rect 13960 19560 14050 19800
rect 14290 19560 14380 19800
rect 14620 19560 14710 19800
rect 14950 19560 15040 19800
rect 15280 19560 15370 19800
rect 15610 19560 15700 19800
rect 15940 19560 16030 19800
rect 16270 19560 16360 19800
rect 16600 19560 16690 19800
rect 16930 19560 17020 19800
rect 17260 19560 17350 19800
rect 17590 19560 17680 19800
rect 17920 19560 18010 19800
rect 18250 19560 18340 19800
rect 18580 19560 18670 19800
rect 18910 19560 19000 19800
rect 19240 19560 19330 19800
rect 19570 19560 19920 19800
rect 7610 19470 19920 19560
rect 7610 19230 7780 19470
rect 8020 19230 8110 19470
rect 8350 19230 8440 19470
rect 8680 19230 8770 19470
rect 9010 19230 9100 19470
rect 9340 19230 9430 19470
rect 9670 19230 9760 19470
rect 10000 19230 10090 19470
rect 10330 19230 10420 19470
rect 10660 19230 10750 19470
rect 10990 19230 11080 19470
rect 11320 19230 11410 19470
rect 11650 19230 11740 19470
rect 11980 19230 12070 19470
rect 12310 19230 12400 19470
rect 12640 19230 12730 19470
rect 12970 19230 13060 19470
rect 13300 19230 13390 19470
rect 13630 19230 13720 19470
rect 13960 19230 14050 19470
rect 14290 19230 14380 19470
rect 14620 19230 14710 19470
rect 14950 19230 15040 19470
rect 15280 19230 15370 19470
rect 15610 19230 15700 19470
rect 15940 19230 16030 19470
rect 16270 19230 16360 19470
rect 16600 19230 16690 19470
rect 16930 19230 17020 19470
rect 17260 19230 17350 19470
rect 17590 19230 17680 19470
rect 17920 19230 18010 19470
rect 18250 19230 18340 19470
rect 18580 19230 18670 19470
rect 18910 19230 19000 19470
rect 19240 19230 19330 19470
rect 19570 19230 19920 19470
rect 7610 19140 19920 19230
rect 7610 18900 7780 19140
rect 8020 18900 8110 19140
rect 8350 18900 8440 19140
rect 8680 18900 8770 19140
rect 9010 18900 9100 19140
rect 9340 18900 9430 19140
rect 9670 18900 9760 19140
rect 10000 18900 10090 19140
rect 10330 18900 10420 19140
rect 10660 18900 10750 19140
rect 10990 18900 11080 19140
rect 11320 18900 11410 19140
rect 11650 18900 11740 19140
rect 11980 18900 12070 19140
rect 12310 18900 12400 19140
rect 12640 18900 12730 19140
rect 12970 18900 13060 19140
rect 13300 18900 13390 19140
rect 13630 18900 13720 19140
rect 13960 18900 14050 19140
rect 14290 18900 14380 19140
rect 14620 18900 14710 19140
rect 14950 18900 15040 19140
rect 15280 18900 15370 19140
rect 15610 18900 15700 19140
rect 15940 18900 16030 19140
rect 16270 18900 16360 19140
rect 16600 18900 16690 19140
rect 16930 18900 17020 19140
rect 17260 18900 17350 19140
rect 17590 18900 17680 19140
rect 17920 18900 18010 19140
rect 18250 18900 18340 19140
rect 18580 18900 18670 19140
rect 18910 18900 19000 19140
rect 19240 18900 19330 19140
rect 19570 18900 19920 19140
rect 7610 18810 19920 18900
rect 7610 18570 7780 18810
rect 8020 18570 8110 18810
rect 8350 18570 8440 18810
rect 8680 18570 8770 18810
rect 9010 18570 9100 18810
rect 9340 18570 9430 18810
rect 9670 18570 9760 18810
rect 10000 18570 10090 18810
rect 10330 18570 10420 18810
rect 10660 18570 10750 18810
rect 10990 18570 11080 18810
rect 11320 18570 11410 18810
rect 11650 18570 11740 18810
rect 11980 18570 12070 18810
rect 12310 18570 12400 18810
rect 12640 18570 12730 18810
rect 12970 18570 13060 18810
rect 13300 18570 13390 18810
rect 13630 18570 13720 18810
rect 13960 18570 14050 18810
rect 14290 18570 14380 18810
rect 14620 18570 14710 18810
rect 14950 18570 15040 18810
rect 15280 18570 15370 18810
rect 15610 18570 15700 18810
rect 15940 18570 16030 18810
rect 16270 18570 16360 18810
rect 16600 18570 16690 18810
rect 16930 18570 17020 18810
rect 17260 18570 17350 18810
rect 17590 18570 17680 18810
rect 17920 18570 18010 18810
rect 18250 18570 18340 18810
rect 18580 18570 18670 18810
rect 18910 18570 19000 18810
rect 19240 18570 19330 18810
rect 19570 18570 19920 18810
rect 7610 18480 19920 18570
rect 7610 18240 7780 18480
rect 8020 18240 8110 18480
rect 8350 18240 8440 18480
rect 8680 18240 8770 18480
rect 9010 18240 9100 18480
rect 9340 18240 9430 18480
rect 9670 18240 9760 18480
rect 10000 18240 10090 18480
rect 10330 18240 10420 18480
rect 10660 18240 10750 18480
rect 10990 18240 11080 18480
rect 11320 18240 11410 18480
rect 11650 18240 11740 18480
rect 11980 18240 12070 18480
rect 12310 18240 12400 18480
rect 12640 18240 12730 18480
rect 12970 18240 13060 18480
rect 13300 18240 13390 18480
rect 13630 18240 13720 18480
rect 13960 18240 14050 18480
rect 14290 18240 14380 18480
rect 14620 18240 14710 18480
rect 14950 18240 15040 18480
rect 15280 18240 15370 18480
rect 15610 18240 15700 18480
rect 15940 18240 16030 18480
rect 16270 18240 16360 18480
rect 16600 18240 16690 18480
rect 16930 18240 17020 18480
rect 17260 18240 17350 18480
rect 17590 18240 17680 18480
rect 17920 18240 18010 18480
rect 18250 18240 18340 18480
rect 18580 18240 18670 18480
rect 18910 18240 19000 18480
rect 19240 18240 19330 18480
rect 19570 18240 19920 18480
rect 7610 18150 19920 18240
rect 7610 17910 7780 18150
rect 8020 17910 8110 18150
rect 8350 17910 8440 18150
rect 8680 17910 8770 18150
rect 9010 17910 9100 18150
rect 9340 17910 9430 18150
rect 9670 17910 9760 18150
rect 10000 17910 10090 18150
rect 10330 17910 10420 18150
rect 10660 17910 10750 18150
rect 10990 17910 11080 18150
rect 11320 17910 11410 18150
rect 11650 17910 11740 18150
rect 11980 17910 12070 18150
rect 12310 17910 12400 18150
rect 12640 17910 12730 18150
rect 12970 17910 13060 18150
rect 13300 17910 13390 18150
rect 13630 17910 13720 18150
rect 13960 17910 14050 18150
rect 14290 17910 14380 18150
rect 14620 17910 14710 18150
rect 14950 17910 15040 18150
rect 15280 17910 15370 18150
rect 15610 17910 15700 18150
rect 15940 17910 16030 18150
rect 16270 17910 16360 18150
rect 16600 17910 16690 18150
rect 16930 17910 17020 18150
rect 17260 17910 17350 18150
rect 17590 17910 17680 18150
rect 17920 17910 18010 18150
rect 18250 17910 18340 18150
rect 18580 17910 18670 18150
rect 18910 17910 19000 18150
rect 19240 17910 19330 18150
rect 19570 17910 19920 18150
rect 7610 17820 19920 17910
rect 7610 17580 7780 17820
rect 8020 17580 8110 17820
rect 8350 17580 8440 17820
rect 8680 17580 8770 17820
rect 9010 17580 9100 17820
rect 9340 17580 9430 17820
rect 9670 17580 9760 17820
rect 10000 17580 10090 17820
rect 10330 17580 10420 17820
rect 10660 17580 10750 17820
rect 10990 17580 11080 17820
rect 11320 17580 11410 17820
rect 11650 17580 11740 17820
rect 11980 17580 12070 17820
rect 12310 17580 12400 17820
rect 12640 17580 12730 17820
rect 12970 17580 13060 17820
rect 13300 17580 13390 17820
rect 13630 17580 13720 17820
rect 13960 17580 14050 17820
rect 14290 17580 14380 17820
rect 14620 17580 14710 17820
rect 14950 17580 15040 17820
rect 15280 17580 15370 17820
rect 15610 17580 15700 17820
rect 15940 17580 16030 17820
rect 16270 17580 16360 17820
rect 16600 17580 16690 17820
rect 16930 17580 17020 17820
rect 17260 17580 17350 17820
rect 17590 17580 17680 17820
rect 17920 17580 18010 17820
rect 18250 17580 18340 17820
rect 18580 17580 18670 17820
rect 18910 17580 19000 17820
rect 19240 17580 19330 17820
rect 19570 17580 19920 17820
rect 7610 17490 19920 17580
rect 7610 17250 7780 17490
rect 8020 17250 8110 17490
rect 8350 17250 8440 17490
rect 8680 17250 8770 17490
rect 9010 17250 9100 17490
rect 9340 17250 9430 17490
rect 9670 17250 9760 17490
rect 10000 17250 10090 17490
rect 10330 17250 10420 17490
rect 10660 17250 10750 17490
rect 10990 17250 11080 17490
rect 11320 17250 11410 17490
rect 11650 17250 11740 17490
rect 11980 17250 12070 17490
rect 12310 17250 12400 17490
rect 12640 17250 12730 17490
rect 12970 17250 13060 17490
rect 13300 17250 13390 17490
rect 13630 17250 13720 17490
rect 13960 17250 14050 17490
rect 14290 17250 14380 17490
rect 14620 17250 14710 17490
rect 14950 17250 15040 17490
rect 15280 17250 15370 17490
rect 15610 17250 15700 17490
rect 15940 17250 16030 17490
rect 16270 17250 16360 17490
rect 16600 17250 16690 17490
rect 16930 17250 17020 17490
rect 17260 17250 17350 17490
rect 17590 17250 17680 17490
rect 17920 17250 18010 17490
rect 18250 17250 18340 17490
rect 18580 17250 18670 17490
rect 18910 17250 19000 17490
rect 19240 17250 19330 17490
rect 19570 17250 19920 17490
rect 7610 17160 19920 17250
rect 7610 16920 7780 17160
rect 8020 16920 8110 17160
rect 8350 16920 8440 17160
rect 8680 16920 8770 17160
rect 9010 16920 9100 17160
rect 9340 16920 9430 17160
rect 9670 16920 9760 17160
rect 10000 16920 10090 17160
rect 10330 16920 10420 17160
rect 10660 16920 10750 17160
rect 10990 16920 11080 17160
rect 11320 16920 11410 17160
rect 11650 16920 11740 17160
rect 11980 16920 12070 17160
rect 12310 16920 12400 17160
rect 12640 16920 12730 17160
rect 12970 16920 13060 17160
rect 13300 16920 13390 17160
rect 13630 16920 13720 17160
rect 13960 16920 14050 17160
rect 14290 16920 14380 17160
rect 14620 16920 14710 17160
rect 14950 16920 15040 17160
rect 15280 16920 15370 17160
rect 15610 16920 15700 17160
rect 15940 16920 16030 17160
rect 16270 16920 16360 17160
rect 16600 16920 16690 17160
rect 16930 16920 17020 17160
rect 17260 16920 17350 17160
rect 17590 16920 17680 17160
rect 17920 16920 18010 17160
rect 18250 16920 18340 17160
rect 18580 16920 18670 17160
rect 18910 16920 19000 17160
rect 19240 16920 19330 17160
rect 19570 16920 19920 17160
rect 7610 16830 19920 16920
rect 7610 16590 7780 16830
rect 8020 16590 8110 16830
rect 8350 16590 8440 16830
rect 8680 16590 8770 16830
rect 9010 16590 9100 16830
rect 9340 16590 9430 16830
rect 9670 16590 9760 16830
rect 10000 16590 10090 16830
rect 10330 16590 10420 16830
rect 10660 16590 10750 16830
rect 10990 16590 11080 16830
rect 11320 16590 11410 16830
rect 11650 16590 11740 16830
rect 11980 16590 12070 16830
rect 12310 16590 12400 16830
rect 12640 16590 12730 16830
rect 12970 16590 13060 16830
rect 13300 16590 13390 16830
rect 13630 16590 13720 16830
rect 13960 16590 14050 16830
rect 14290 16590 14380 16830
rect 14620 16590 14710 16830
rect 14950 16590 15040 16830
rect 15280 16590 15370 16830
rect 15610 16590 15700 16830
rect 15940 16590 16030 16830
rect 16270 16590 16360 16830
rect 16600 16590 16690 16830
rect 16930 16590 17020 16830
rect 17260 16590 17350 16830
rect 17590 16590 17680 16830
rect 17920 16590 18010 16830
rect 18250 16590 18340 16830
rect 18580 16590 18670 16830
rect 18910 16590 19000 16830
rect 19240 16590 19330 16830
rect 19570 16590 19920 16830
rect 7610 16500 19920 16590
rect 7610 16260 7780 16500
rect 8020 16260 8110 16500
rect 8350 16260 8440 16500
rect 8680 16260 8770 16500
rect 9010 16260 9100 16500
rect 9340 16260 9430 16500
rect 9670 16260 9760 16500
rect 10000 16260 10090 16500
rect 10330 16260 10420 16500
rect 10660 16260 10750 16500
rect 10990 16260 11080 16500
rect 11320 16260 11410 16500
rect 11650 16260 11740 16500
rect 11980 16260 12070 16500
rect 12310 16260 12400 16500
rect 12640 16260 12730 16500
rect 12970 16260 13060 16500
rect 13300 16260 13390 16500
rect 13630 16260 13720 16500
rect 13960 16260 14050 16500
rect 14290 16260 14380 16500
rect 14620 16260 14710 16500
rect 14950 16260 15040 16500
rect 15280 16260 15370 16500
rect 15610 16260 15700 16500
rect 15940 16260 16030 16500
rect 16270 16260 16360 16500
rect 16600 16260 16690 16500
rect 16930 16260 17020 16500
rect 17260 16260 17350 16500
rect 17590 16260 17680 16500
rect 17920 16260 18010 16500
rect 18250 16260 18340 16500
rect 18580 16260 18670 16500
rect 18910 16260 19000 16500
rect 19240 16260 19330 16500
rect 19570 16260 19920 16500
rect 7610 16170 19920 16260
rect 7610 15930 7780 16170
rect 8020 15930 8110 16170
rect 8350 15930 8440 16170
rect 8680 15930 8770 16170
rect 9010 15930 9100 16170
rect 9340 15930 9430 16170
rect 9670 15930 9760 16170
rect 10000 15930 10090 16170
rect 10330 15930 10420 16170
rect 10660 15930 10750 16170
rect 10990 15930 11080 16170
rect 11320 15930 11410 16170
rect 11650 15930 11740 16170
rect 11980 15930 12070 16170
rect 12310 15930 12400 16170
rect 12640 15930 12730 16170
rect 12970 15930 13060 16170
rect 13300 15930 13390 16170
rect 13630 15930 13720 16170
rect 13960 15930 14050 16170
rect 14290 15930 14380 16170
rect 14620 15930 14710 16170
rect 14950 15930 15040 16170
rect 15280 15930 15370 16170
rect 15610 15930 15700 16170
rect 15940 15930 16030 16170
rect 16270 15930 16360 16170
rect 16600 15930 16690 16170
rect 16930 15930 17020 16170
rect 17260 15930 17350 16170
rect 17590 15930 17680 16170
rect 17920 15930 18010 16170
rect 18250 15930 18340 16170
rect 18580 15930 18670 16170
rect 18910 15930 19000 16170
rect 19240 15930 19330 16170
rect 19570 15930 19920 16170
rect 7610 15840 19920 15930
rect 7610 15600 7780 15840
rect 8020 15600 8110 15840
rect 8350 15600 8440 15840
rect 8680 15600 8770 15840
rect 9010 15600 9100 15840
rect 9340 15600 9430 15840
rect 9670 15600 9760 15840
rect 10000 15600 10090 15840
rect 10330 15600 10420 15840
rect 10660 15600 10750 15840
rect 10990 15600 11080 15840
rect 11320 15600 11410 15840
rect 11650 15600 11740 15840
rect 11980 15600 12070 15840
rect 12310 15600 12400 15840
rect 12640 15600 12730 15840
rect 12970 15600 13060 15840
rect 13300 15600 13390 15840
rect 13630 15600 13720 15840
rect 13960 15600 14050 15840
rect 14290 15600 14380 15840
rect 14620 15600 14710 15840
rect 14950 15600 15040 15840
rect 15280 15600 15370 15840
rect 15610 15600 15700 15840
rect 15940 15600 16030 15840
rect 16270 15600 16360 15840
rect 16600 15600 16690 15840
rect 16930 15600 17020 15840
rect 17260 15600 17350 15840
rect 17590 15600 17680 15840
rect 17920 15600 18010 15840
rect 18250 15600 18340 15840
rect 18580 15600 18670 15840
rect 18910 15600 19000 15840
rect 19240 15600 19330 15840
rect 19570 15600 19920 15840
rect 7610 15510 19920 15600
rect 7610 15270 7780 15510
rect 8020 15270 8110 15510
rect 8350 15270 8440 15510
rect 8680 15270 8770 15510
rect 9010 15270 9100 15510
rect 9340 15270 9430 15510
rect 9670 15270 9760 15510
rect 10000 15270 10090 15510
rect 10330 15270 10420 15510
rect 10660 15270 10750 15510
rect 10990 15270 11080 15510
rect 11320 15270 11410 15510
rect 11650 15270 11740 15510
rect 11980 15270 12070 15510
rect 12310 15270 12400 15510
rect 12640 15270 12730 15510
rect 12970 15270 13060 15510
rect 13300 15270 13390 15510
rect 13630 15270 13720 15510
rect 13960 15270 14050 15510
rect 14290 15270 14380 15510
rect 14620 15270 14710 15510
rect 14950 15270 15040 15510
rect 15280 15270 15370 15510
rect 15610 15270 15700 15510
rect 15940 15270 16030 15510
rect 16270 15270 16360 15510
rect 16600 15270 16690 15510
rect 16930 15270 17020 15510
rect 17260 15270 17350 15510
rect 17590 15270 17680 15510
rect 17920 15270 18010 15510
rect 18250 15270 18340 15510
rect 18580 15270 18670 15510
rect 18910 15270 19000 15510
rect 19240 15270 19330 15510
rect 19570 15270 19920 15510
rect 7610 15180 19920 15270
rect 7610 14940 7780 15180
rect 8020 14940 8110 15180
rect 8350 14940 8440 15180
rect 8680 14940 8770 15180
rect 9010 14940 9100 15180
rect 9340 14940 9430 15180
rect 9670 14940 9760 15180
rect 10000 14940 10090 15180
rect 10330 14940 10420 15180
rect 10660 14940 10750 15180
rect 10990 14940 11080 15180
rect 11320 14940 11410 15180
rect 11650 14940 11740 15180
rect 11980 14940 12070 15180
rect 12310 14940 12400 15180
rect 12640 14940 12730 15180
rect 12970 14940 13060 15180
rect 13300 14940 13390 15180
rect 13630 14940 13720 15180
rect 13960 14940 14050 15180
rect 14290 14940 14380 15180
rect 14620 14940 14710 15180
rect 14950 14940 15040 15180
rect 15280 14940 15370 15180
rect 15610 14940 15700 15180
rect 15940 14940 16030 15180
rect 16270 14940 16360 15180
rect 16600 14940 16690 15180
rect 16930 14940 17020 15180
rect 17260 14940 17350 15180
rect 17590 14940 17680 15180
rect 17920 14940 18010 15180
rect 18250 14940 18340 15180
rect 18580 14940 18670 15180
rect 18910 14940 19000 15180
rect 19240 14940 19330 15180
rect 19570 14940 19920 15180
rect 7610 14850 19920 14940
rect 7610 14610 7780 14850
rect 8020 14610 8110 14850
rect 8350 14610 8440 14850
rect 8680 14610 8770 14850
rect 9010 14610 9100 14850
rect 9340 14610 9430 14850
rect 9670 14610 9760 14850
rect 10000 14610 10090 14850
rect 10330 14610 10420 14850
rect 10660 14610 10750 14850
rect 10990 14610 11080 14850
rect 11320 14610 11410 14850
rect 11650 14610 11740 14850
rect 11980 14610 12070 14850
rect 12310 14610 12400 14850
rect 12640 14610 12730 14850
rect 12970 14610 13060 14850
rect 13300 14610 13390 14850
rect 13630 14610 13720 14850
rect 13960 14610 14050 14850
rect 14290 14610 14380 14850
rect 14620 14610 14710 14850
rect 14950 14610 15040 14850
rect 15280 14610 15370 14850
rect 15610 14610 15700 14850
rect 15940 14610 16030 14850
rect 16270 14610 16360 14850
rect 16600 14610 16690 14850
rect 16930 14610 17020 14850
rect 17260 14610 17350 14850
rect 17590 14610 17680 14850
rect 17920 14610 18010 14850
rect 18250 14610 18340 14850
rect 18580 14610 18670 14850
rect 18910 14610 19000 14850
rect 19240 14610 19330 14850
rect 19570 14610 19920 14850
rect 7610 14520 19920 14610
rect 7610 14280 7780 14520
rect 8020 14280 8110 14520
rect 8350 14280 8440 14520
rect 8680 14280 8770 14520
rect 9010 14280 9100 14520
rect 9340 14280 9430 14520
rect 9670 14280 9760 14520
rect 10000 14280 10090 14520
rect 10330 14280 10420 14520
rect 10660 14280 10750 14520
rect 10990 14280 11080 14520
rect 11320 14280 11410 14520
rect 11650 14280 11740 14520
rect 11980 14280 12070 14520
rect 12310 14280 12400 14520
rect 12640 14280 12730 14520
rect 12970 14280 13060 14520
rect 13300 14280 13390 14520
rect 13630 14280 13720 14520
rect 13960 14280 14050 14520
rect 14290 14280 14380 14520
rect 14620 14280 14710 14520
rect 14950 14280 15040 14520
rect 15280 14280 15370 14520
rect 15610 14280 15700 14520
rect 15940 14280 16030 14520
rect 16270 14280 16360 14520
rect 16600 14280 16690 14520
rect 16930 14280 17020 14520
rect 17260 14280 17350 14520
rect 17590 14280 17680 14520
rect 17920 14280 18010 14520
rect 18250 14280 18340 14520
rect 18580 14280 18670 14520
rect 18910 14280 19000 14520
rect 19240 14280 19330 14520
rect 19570 14280 19920 14520
rect 7610 14190 19920 14280
rect 7610 13950 7780 14190
rect 8020 13950 8110 14190
rect 8350 13950 8440 14190
rect 8680 13950 8770 14190
rect 9010 13950 9100 14190
rect 9340 13950 9430 14190
rect 9670 13950 9760 14190
rect 10000 13950 10090 14190
rect 10330 13950 10420 14190
rect 10660 13950 10750 14190
rect 10990 13950 11080 14190
rect 11320 13950 11410 14190
rect 11650 13950 11740 14190
rect 11980 13950 12070 14190
rect 12310 13950 12400 14190
rect 12640 13950 12730 14190
rect 12970 13950 13060 14190
rect 13300 13950 13390 14190
rect 13630 13950 13720 14190
rect 13960 13950 14050 14190
rect 14290 13950 14380 14190
rect 14620 13950 14710 14190
rect 14950 13950 15040 14190
rect 15280 13950 15370 14190
rect 15610 13950 15700 14190
rect 15940 13950 16030 14190
rect 16270 13950 16360 14190
rect 16600 13950 16690 14190
rect 16930 13950 17020 14190
rect 17260 13950 17350 14190
rect 17590 13950 17680 14190
rect 17920 13950 18010 14190
rect 18250 13950 18340 14190
rect 18580 13950 18670 14190
rect 18910 13950 19000 14190
rect 19240 13950 19330 14190
rect 19570 13950 19920 14190
rect 7610 13860 19920 13950
rect 7610 13620 7780 13860
rect 8020 13620 8110 13860
rect 8350 13620 8440 13860
rect 8680 13620 8770 13860
rect 9010 13620 9100 13860
rect 9340 13620 9430 13860
rect 9670 13620 9760 13860
rect 10000 13620 10090 13860
rect 10330 13620 10420 13860
rect 10660 13620 10750 13860
rect 10990 13620 11080 13860
rect 11320 13620 11410 13860
rect 11650 13620 11740 13860
rect 11980 13620 12070 13860
rect 12310 13620 12400 13860
rect 12640 13620 12730 13860
rect 12970 13620 13060 13860
rect 13300 13620 13390 13860
rect 13630 13620 13720 13860
rect 13960 13620 14050 13860
rect 14290 13620 14380 13860
rect 14620 13620 14710 13860
rect 14950 13620 15040 13860
rect 15280 13620 15370 13860
rect 15610 13620 15700 13860
rect 15940 13620 16030 13860
rect 16270 13620 16360 13860
rect 16600 13620 16690 13860
rect 16930 13620 17020 13860
rect 17260 13620 17350 13860
rect 17590 13620 17680 13860
rect 17920 13620 18010 13860
rect 18250 13620 18340 13860
rect 18580 13620 18670 13860
rect 18910 13620 19000 13860
rect 19240 13620 19330 13860
rect 19570 13620 19920 13860
rect 7610 13530 19920 13620
rect 7610 13290 7780 13530
rect 8020 13290 8110 13530
rect 8350 13290 8440 13530
rect 8680 13290 8770 13530
rect 9010 13290 9100 13530
rect 9340 13290 9430 13530
rect 9670 13290 9760 13530
rect 10000 13290 10090 13530
rect 10330 13290 10420 13530
rect 10660 13290 10750 13530
rect 10990 13290 11080 13530
rect 11320 13290 11410 13530
rect 11650 13290 11740 13530
rect 11980 13290 12070 13530
rect 12310 13290 12400 13530
rect 12640 13290 12730 13530
rect 12970 13290 13060 13530
rect 13300 13290 13390 13530
rect 13630 13290 13720 13530
rect 13960 13290 14050 13530
rect 14290 13290 14380 13530
rect 14620 13290 14710 13530
rect 14950 13290 15040 13530
rect 15280 13290 15370 13530
rect 15610 13290 15700 13530
rect 15940 13290 16030 13530
rect 16270 13290 16360 13530
rect 16600 13290 16690 13530
rect 16930 13290 17020 13530
rect 17260 13290 17350 13530
rect 17590 13290 17680 13530
rect 17920 13290 18010 13530
rect 18250 13290 18340 13530
rect 18580 13290 18670 13530
rect 18910 13290 19000 13530
rect 19240 13290 19330 13530
rect 19570 13290 19920 13530
rect 7610 13200 19920 13290
rect 7610 12960 7780 13200
rect 8020 12960 8110 13200
rect 8350 12960 8440 13200
rect 8680 12960 8770 13200
rect 9010 12960 9100 13200
rect 9340 12960 9430 13200
rect 9670 12960 9760 13200
rect 10000 12960 10090 13200
rect 10330 12960 10420 13200
rect 10660 12960 10750 13200
rect 10990 12960 11080 13200
rect 11320 12960 11410 13200
rect 11650 12960 11740 13200
rect 11980 12960 12070 13200
rect 12310 12960 12400 13200
rect 12640 12960 12730 13200
rect 12970 12960 13060 13200
rect 13300 12960 13390 13200
rect 13630 12960 13720 13200
rect 13960 12960 14050 13200
rect 14290 12960 14380 13200
rect 14620 12960 14710 13200
rect 14950 12960 15040 13200
rect 15280 12960 15370 13200
rect 15610 12960 15700 13200
rect 15940 12960 16030 13200
rect 16270 12960 16360 13200
rect 16600 12960 16690 13200
rect 16930 12960 17020 13200
rect 17260 12960 17350 13200
rect 17590 12960 17680 13200
rect 17920 12960 18010 13200
rect 18250 12960 18340 13200
rect 18580 12960 18670 13200
rect 18910 12960 19000 13200
rect 19240 12960 19330 13200
rect 19570 12960 19920 13200
rect 7610 12870 19920 12960
rect 7610 12630 7780 12870
rect 8020 12630 8110 12870
rect 8350 12630 8440 12870
rect 8680 12630 8770 12870
rect 9010 12630 9100 12870
rect 9340 12630 9430 12870
rect 9670 12630 9760 12870
rect 10000 12630 10090 12870
rect 10330 12630 10420 12870
rect 10660 12630 10750 12870
rect 10990 12630 11080 12870
rect 11320 12630 11410 12870
rect 11650 12630 11740 12870
rect 11980 12630 12070 12870
rect 12310 12630 12400 12870
rect 12640 12630 12730 12870
rect 12970 12630 13060 12870
rect 13300 12630 13390 12870
rect 13630 12630 13720 12870
rect 13960 12630 14050 12870
rect 14290 12630 14380 12870
rect 14620 12630 14710 12870
rect 14950 12630 15040 12870
rect 15280 12630 15370 12870
rect 15610 12630 15700 12870
rect 15940 12630 16030 12870
rect 16270 12630 16360 12870
rect 16600 12630 16690 12870
rect 16930 12630 17020 12870
rect 17260 12630 17350 12870
rect 17590 12630 17680 12870
rect 17920 12630 18010 12870
rect 18250 12630 18340 12870
rect 18580 12630 18670 12870
rect 18910 12630 19000 12870
rect 19240 12630 19330 12870
rect 19570 12630 19920 12870
rect 7610 12540 19920 12630
rect 7610 12300 7780 12540
rect 8020 12300 8110 12540
rect 8350 12300 8440 12540
rect 8680 12300 8770 12540
rect 9010 12300 9100 12540
rect 9340 12300 9430 12540
rect 9670 12300 9760 12540
rect 10000 12300 10090 12540
rect 10330 12300 10420 12540
rect 10660 12300 10750 12540
rect 10990 12300 11080 12540
rect 11320 12300 11410 12540
rect 11650 12300 11740 12540
rect 11980 12300 12070 12540
rect 12310 12300 12400 12540
rect 12640 12300 12730 12540
rect 12970 12300 13060 12540
rect 13300 12300 13390 12540
rect 13630 12300 13720 12540
rect 13960 12300 14050 12540
rect 14290 12300 14380 12540
rect 14620 12300 14710 12540
rect 14950 12300 15040 12540
rect 15280 12300 15370 12540
rect 15610 12300 15700 12540
rect 15940 12300 16030 12540
rect 16270 12300 16360 12540
rect 16600 12300 16690 12540
rect 16930 12300 17020 12540
rect 17260 12300 17350 12540
rect 17590 12300 17680 12540
rect 17920 12300 18010 12540
rect 18250 12300 18340 12540
rect 18580 12300 18670 12540
rect 18910 12300 19000 12540
rect 19240 12300 19330 12540
rect 19570 12300 19920 12540
rect 7610 12210 19920 12300
rect 7610 11970 7780 12210
rect 8020 11970 8110 12210
rect 8350 11970 8440 12210
rect 8680 11970 8770 12210
rect 9010 11970 9100 12210
rect 9340 11970 9430 12210
rect 9670 11970 9760 12210
rect 10000 11970 10090 12210
rect 10330 11970 10420 12210
rect 10660 11970 10750 12210
rect 10990 11970 11080 12210
rect 11320 11970 11410 12210
rect 11650 11970 11740 12210
rect 11980 11970 12070 12210
rect 12310 11970 12400 12210
rect 12640 11970 12730 12210
rect 12970 11970 13060 12210
rect 13300 11970 13390 12210
rect 13630 11970 13720 12210
rect 13960 11970 14050 12210
rect 14290 11970 14380 12210
rect 14620 11970 14710 12210
rect 14950 11970 15040 12210
rect 15280 11970 15370 12210
rect 15610 11970 15700 12210
rect 15940 11970 16030 12210
rect 16270 11970 16360 12210
rect 16600 11970 16690 12210
rect 16930 11970 17020 12210
rect 17260 11970 17350 12210
rect 17590 11970 17680 12210
rect 17920 11970 18010 12210
rect 18250 11970 18340 12210
rect 18580 11970 18670 12210
rect 18910 11970 19000 12210
rect 19240 11970 19330 12210
rect 19570 11970 19920 12210
rect 7610 11880 19920 11970
rect 7610 11640 7780 11880
rect 8020 11640 8110 11880
rect 8350 11640 8440 11880
rect 8680 11640 8770 11880
rect 9010 11640 9100 11880
rect 9340 11640 9430 11880
rect 9670 11640 9760 11880
rect 10000 11640 10090 11880
rect 10330 11640 10420 11880
rect 10660 11640 10750 11880
rect 10990 11640 11080 11880
rect 11320 11640 11410 11880
rect 11650 11640 11740 11880
rect 11980 11640 12070 11880
rect 12310 11640 12400 11880
rect 12640 11640 12730 11880
rect 12970 11640 13060 11880
rect 13300 11640 13390 11880
rect 13630 11640 13720 11880
rect 13960 11640 14050 11880
rect 14290 11640 14380 11880
rect 14620 11640 14710 11880
rect 14950 11640 15040 11880
rect 15280 11640 15370 11880
rect 15610 11640 15700 11880
rect 15940 11640 16030 11880
rect 16270 11640 16360 11880
rect 16600 11640 16690 11880
rect 16930 11640 17020 11880
rect 17260 11640 17350 11880
rect 17590 11640 17680 11880
rect 17920 11640 18010 11880
rect 18250 11640 18340 11880
rect 18580 11640 18670 11880
rect 18910 11640 19000 11880
rect 19240 11640 19330 11880
rect 19570 11640 19920 11880
rect 7610 11550 19920 11640
rect 7610 11310 7780 11550
rect 8020 11310 8110 11550
rect 8350 11310 8440 11550
rect 8680 11310 8770 11550
rect 9010 11310 9100 11550
rect 9340 11310 9430 11550
rect 9670 11310 9760 11550
rect 10000 11310 10090 11550
rect 10330 11310 10420 11550
rect 10660 11310 10750 11550
rect 10990 11310 11080 11550
rect 11320 11310 11410 11550
rect 11650 11310 11740 11550
rect 11980 11310 12070 11550
rect 12310 11310 12400 11550
rect 12640 11310 12730 11550
rect 12970 11310 13060 11550
rect 13300 11310 13390 11550
rect 13630 11310 13720 11550
rect 13960 11310 14050 11550
rect 14290 11310 14380 11550
rect 14620 11310 14710 11550
rect 14950 11310 15040 11550
rect 15280 11310 15370 11550
rect 15610 11310 15700 11550
rect 15940 11310 16030 11550
rect 16270 11310 16360 11550
rect 16600 11310 16690 11550
rect 16930 11310 17020 11550
rect 17260 11310 17350 11550
rect 17590 11310 17680 11550
rect 17920 11310 18010 11550
rect 18250 11310 18340 11550
rect 18580 11310 18670 11550
rect 18910 11310 19000 11550
rect 19240 11310 19330 11550
rect 19570 11310 19920 11550
rect 7610 11220 19920 11310
rect 7610 10980 7780 11220
rect 8020 10980 8110 11220
rect 8350 10980 8440 11220
rect 8680 10980 8770 11220
rect 9010 10980 9100 11220
rect 9340 10980 9430 11220
rect 9670 10980 9760 11220
rect 10000 10980 10090 11220
rect 10330 10980 10420 11220
rect 10660 10980 10750 11220
rect 10990 10980 11080 11220
rect 11320 10980 11410 11220
rect 11650 10980 11740 11220
rect 11980 10980 12070 11220
rect 12310 10980 12400 11220
rect 12640 10980 12730 11220
rect 12970 10980 13060 11220
rect 13300 10980 13390 11220
rect 13630 10980 13720 11220
rect 13960 10980 14050 11220
rect 14290 10980 14380 11220
rect 14620 10980 14710 11220
rect 14950 10980 15040 11220
rect 15280 10980 15370 11220
rect 15610 10980 15700 11220
rect 15940 10980 16030 11220
rect 16270 10980 16360 11220
rect 16600 10980 16690 11220
rect 16930 10980 17020 11220
rect 17260 10980 17350 11220
rect 17590 10980 17680 11220
rect 17920 10980 18010 11220
rect 18250 10980 18340 11220
rect 18580 10980 18670 11220
rect 18910 10980 19000 11220
rect 19240 10980 19330 11220
rect 19570 10980 19920 11220
rect 7610 10890 19920 10980
rect 7610 10650 7780 10890
rect 8020 10650 8110 10890
rect 8350 10650 8440 10890
rect 8680 10650 8770 10890
rect 9010 10650 9100 10890
rect 9340 10650 9430 10890
rect 9670 10650 9760 10890
rect 10000 10650 10090 10890
rect 10330 10650 10420 10890
rect 10660 10650 10750 10890
rect 10990 10650 11080 10890
rect 11320 10650 11410 10890
rect 11650 10650 11740 10890
rect 11980 10650 12070 10890
rect 12310 10650 12400 10890
rect 12640 10650 12730 10890
rect 12970 10650 13060 10890
rect 13300 10650 13390 10890
rect 13630 10650 13720 10890
rect 13960 10650 14050 10890
rect 14290 10650 14380 10890
rect 14620 10650 14710 10890
rect 14950 10650 15040 10890
rect 15280 10650 15370 10890
rect 15610 10650 15700 10890
rect 15940 10650 16030 10890
rect 16270 10650 16360 10890
rect 16600 10650 16690 10890
rect 16930 10650 17020 10890
rect 17260 10650 17350 10890
rect 17590 10650 17680 10890
rect 17920 10650 18010 10890
rect 18250 10650 18340 10890
rect 18580 10650 18670 10890
rect 18910 10650 19000 10890
rect 19240 10650 19330 10890
rect 19570 10650 19920 10890
rect 7610 10560 19920 10650
rect 7610 10320 7780 10560
rect 8020 10320 8110 10560
rect 8350 10320 8440 10560
rect 8680 10320 8770 10560
rect 9010 10320 9100 10560
rect 9340 10320 9430 10560
rect 9670 10320 9760 10560
rect 10000 10320 10090 10560
rect 10330 10320 10420 10560
rect 10660 10320 10750 10560
rect 10990 10320 11080 10560
rect 11320 10320 11410 10560
rect 11650 10320 11740 10560
rect 11980 10320 12070 10560
rect 12310 10320 12400 10560
rect 12640 10320 12730 10560
rect 12970 10320 13060 10560
rect 13300 10320 13390 10560
rect 13630 10320 13720 10560
rect 13960 10320 14050 10560
rect 14290 10320 14380 10560
rect 14620 10320 14710 10560
rect 14950 10320 15040 10560
rect 15280 10320 15370 10560
rect 15610 10320 15700 10560
rect 15940 10320 16030 10560
rect 16270 10320 16360 10560
rect 16600 10320 16690 10560
rect 16930 10320 17020 10560
rect 17260 10320 17350 10560
rect 17590 10320 17680 10560
rect 17920 10320 18010 10560
rect 18250 10320 18340 10560
rect 18580 10320 18670 10560
rect 18910 10320 19000 10560
rect 19240 10320 19330 10560
rect 19570 10320 19920 10560
rect 7610 10230 19920 10320
rect 7610 9990 7780 10230
rect 8020 9990 8110 10230
rect 8350 9990 8440 10230
rect 8680 9990 8770 10230
rect 9010 9990 9100 10230
rect 9340 9990 9430 10230
rect 9670 9990 9760 10230
rect 10000 9990 10090 10230
rect 10330 9990 10420 10230
rect 10660 9990 10750 10230
rect 10990 9990 11080 10230
rect 11320 9990 11410 10230
rect 11650 9990 11740 10230
rect 11980 9990 12070 10230
rect 12310 9990 12400 10230
rect 12640 9990 12730 10230
rect 12970 9990 13060 10230
rect 13300 9990 13390 10230
rect 13630 9990 13720 10230
rect 13960 9990 14050 10230
rect 14290 9990 14380 10230
rect 14620 9990 14710 10230
rect 14950 9990 15040 10230
rect 15280 9990 15370 10230
rect 15610 9990 15700 10230
rect 15940 9990 16030 10230
rect 16270 9990 16360 10230
rect 16600 9990 16690 10230
rect 16930 9990 17020 10230
rect 17260 9990 17350 10230
rect 17590 9990 17680 10230
rect 17920 9990 18010 10230
rect 18250 9990 18340 10230
rect 18580 9990 18670 10230
rect 18910 9990 19000 10230
rect 19240 9990 19330 10230
rect 19570 9990 19920 10230
rect 7610 9900 19920 9990
rect 7610 9660 7780 9900
rect 8020 9660 8110 9900
rect 8350 9660 8440 9900
rect 8680 9660 8770 9900
rect 9010 9660 9100 9900
rect 9340 9660 9430 9900
rect 9670 9660 9760 9900
rect 10000 9660 10090 9900
rect 10330 9660 10420 9900
rect 10660 9660 10750 9900
rect 10990 9660 11080 9900
rect 11320 9660 11410 9900
rect 11650 9660 11740 9900
rect 11980 9660 12070 9900
rect 12310 9660 12400 9900
rect 12640 9660 12730 9900
rect 12970 9660 13060 9900
rect 13300 9660 13390 9900
rect 13630 9660 13720 9900
rect 13960 9660 14050 9900
rect 14290 9660 14380 9900
rect 14620 9660 14710 9900
rect 14950 9660 15040 9900
rect 15280 9660 15370 9900
rect 15610 9660 15700 9900
rect 15940 9660 16030 9900
rect 16270 9660 16360 9900
rect 16600 9660 16690 9900
rect 16930 9660 17020 9900
rect 17260 9660 17350 9900
rect 17590 9660 17680 9900
rect 17920 9660 18010 9900
rect 18250 9660 18340 9900
rect 18580 9660 18670 9900
rect 18910 9660 19000 9900
rect 19240 9660 19330 9900
rect 19570 9660 19920 9900
rect 7610 9570 19920 9660
rect 7610 9330 7780 9570
rect 8020 9330 8110 9570
rect 8350 9330 8440 9570
rect 8680 9330 8770 9570
rect 9010 9330 9100 9570
rect 9340 9330 9430 9570
rect 9670 9330 9760 9570
rect 10000 9330 10090 9570
rect 10330 9330 10420 9570
rect 10660 9330 10750 9570
rect 10990 9330 11080 9570
rect 11320 9330 11410 9570
rect 11650 9330 11740 9570
rect 11980 9330 12070 9570
rect 12310 9330 12400 9570
rect 12640 9330 12730 9570
rect 12970 9330 13060 9570
rect 13300 9330 13390 9570
rect 13630 9330 13720 9570
rect 13960 9330 14050 9570
rect 14290 9330 14380 9570
rect 14620 9330 14710 9570
rect 14950 9330 15040 9570
rect 15280 9330 15370 9570
rect 15610 9330 15700 9570
rect 15940 9330 16030 9570
rect 16270 9330 16360 9570
rect 16600 9330 16690 9570
rect 16930 9330 17020 9570
rect 17260 9330 17350 9570
rect 17590 9330 17680 9570
rect 17920 9330 18010 9570
rect 18250 9330 18340 9570
rect 18580 9330 18670 9570
rect 18910 9330 19000 9570
rect 19240 9330 19330 9570
rect 19570 9330 19920 9570
rect 7610 9240 19920 9330
rect 7610 9000 7780 9240
rect 8020 9000 8110 9240
rect 8350 9000 8440 9240
rect 8680 9000 8770 9240
rect 9010 9000 9100 9240
rect 9340 9000 9430 9240
rect 9670 9000 9760 9240
rect 10000 9000 10090 9240
rect 10330 9000 10420 9240
rect 10660 9000 10750 9240
rect 10990 9000 11080 9240
rect 11320 9000 11410 9240
rect 11650 9000 11740 9240
rect 11980 9000 12070 9240
rect 12310 9000 12400 9240
rect 12640 9000 12730 9240
rect 12970 9000 13060 9240
rect 13300 9000 13390 9240
rect 13630 9000 13720 9240
rect 13960 9000 14050 9240
rect 14290 9000 14380 9240
rect 14620 9000 14710 9240
rect 14950 9000 15040 9240
rect 15280 9000 15370 9240
rect 15610 9000 15700 9240
rect 15940 9000 16030 9240
rect 16270 9000 16360 9240
rect 16600 9000 16690 9240
rect 16930 9000 17020 9240
rect 17260 9000 17350 9240
rect 17590 9000 17680 9240
rect 17920 9000 18010 9240
rect 18250 9000 18340 9240
rect 18580 9000 18670 9240
rect 18910 9000 19000 9240
rect 19240 9000 19330 9240
rect 19570 9000 19920 9240
rect 7610 8460 19920 9000
rect 7610 8220 7640 8460
rect 7880 8220 7970 8460
rect 8210 8220 8300 8460
rect 8540 8220 8630 8460
rect 8870 8220 8960 8460
rect 9200 8220 9290 8460
rect 9530 8220 9620 8460
rect 9860 8220 9950 8460
rect 10190 8220 10280 8460
rect 10520 8220 10650 8460
rect 10890 8220 10980 8460
rect 11220 8220 11310 8460
rect 11550 8220 11640 8460
rect 11880 8220 11970 8460
rect 12210 8220 12300 8460
rect 12540 8220 12630 8460
rect 12870 8220 12960 8460
rect 13200 8220 13290 8460
rect 13530 8220 13660 8460
rect 13900 8220 13990 8460
rect 14230 8220 14320 8460
rect 14560 8220 14650 8460
rect 14890 8220 14980 8460
rect 15220 8220 15310 8460
rect 15550 8220 15640 8460
rect 15880 8220 15970 8460
rect 16210 8220 16300 8460
rect 16540 8220 16670 8460
rect 16910 8220 17000 8460
rect 17240 8220 17330 8460
rect 17570 8220 17660 8460
rect 17900 8220 17990 8460
rect 18230 8220 18320 8460
rect 18560 8220 18650 8460
rect 18890 8220 18980 8460
rect 19220 8220 19310 8460
rect 19550 8220 19920 8460
rect 7610 8190 19920 8220
rect 28700 7830 36100 7910
rect -6530 6940 14510 7700
rect 28700 7590 28780 7830
rect 29020 7590 29110 7830
rect 29350 7590 29440 7830
rect 29680 7590 29770 7830
rect 30010 7590 30100 7830
rect 30340 7590 30430 7830
rect 30670 7590 30760 7830
rect 31000 7590 31090 7830
rect 31330 7590 31420 7830
rect 31660 7590 31750 7830
rect 31990 7590 32080 7830
rect 32320 7590 32410 7830
rect 32650 7590 32740 7830
rect 32980 7590 33070 7830
rect 33310 7590 33400 7830
rect 33640 7590 33730 7830
rect 33970 7590 34060 7830
rect 34300 7590 34390 7830
rect 34630 7590 34720 7830
rect 34960 7590 35050 7830
rect 35290 7770 36100 7830
rect 35290 7590 35830 7770
rect 28700 7530 35830 7590
rect 36070 7530 36100 7770
rect 28700 7500 36100 7530
rect -6530 6910 11940 6940
rect -6530 6900 1720 6910
rect -6530 -2160 -2530 6900
rect 1540 6670 1720 6900
rect 1960 6670 2050 6910
rect 2290 6670 2390 6910
rect 2630 6670 2720 6910
rect 2960 6900 11940 6910
rect 2960 6670 3140 6900
rect 11760 6700 11940 6900
rect 12180 6700 12270 6940
rect 12510 6700 12610 6940
rect 12850 6700 12940 6940
rect 13180 6900 14510 6940
rect 13180 6700 13360 6900
rect 11760 6670 13360 6700
rect 1540 6640 3140 6670
rect 15210 2500 19210 7310
rect 19570 7270 26870 7500
rect 19570 7100 21110 7270
rect 21060 7030 21110 7100
rect 21480 7100 23510 7270
rect 21480 7030 21540 7100
rect 21060 7000 21540 7030
rect 23460 7030 23510 7100
rect 23880 7100 26870 7270
rect 23880 7030 23940 7100
rect 23460 7000 23940 7030
rect 20020 2600 20500 2630
rect 20020 2500 20080 2600
rect 15210 2360 20080 2500
rect 20450 2500 20500 2600
rect 24500 2600 24980 2630
rect 24500 2500 24560 2600
rect 20450 2360 24560 2500
rect 24930 2360 24980 2600
rect 15210 2100 24980 2360
rect 1080 -790 2680 -760
rect 1080 -1030 1260 -790
rect 1500 -1030 1590 -790
rect 1830 -1030 1930 -790
rect 2170 -1030 2260 -790
rect 2500 -1030 2680 -790
rect 1080 -1040 2680 -1030
rect 12220 -790 13820 -760
rect 12220 -1030 12400 -790
rect 12640 -1030 12730 -790
rect 12970 -1030 13070 -790
rect 13310 -1030 13400 -790
rect 13640 -1030 13820 -790
rect 12220 -1040 13820 -1030
rect 15210 -1040 19210 2100
rect 26180 1440 26870 7100
rect 19680 1040 26870 1440
rect 28700 7260 28780 7500
rect 29020 7260 29110 7500
rect 29350 7260 29440 7500
rect 29680 7260 29770 7500
rect 30010 7260 30100 7500
rect 30340 7260 30430 7500
rect 30670 7260 30760 7500
rect 31000 7260 31090 7500
rect 31330 7260 31420 7500
rect 31660 7260 31750 7500
rect 31990 7260 32080 7500
rect 32320 7260 32410 7500
rect 32650 7260 32740 7500
rect 32980 7260 33070 7500
rect 33310 7260 33400 7500
rect 33640 7260 33730 7500
rect 33970 7260 34060 7500
rect 34300 7260 34390 7500
rect 34630 7260 34720 7500
rect 34960 7260 35050 7500
rect 35290 7440 36100 7500
rect 35290 7260 35830 7440
rect 28700 7200 35830 7260
rect 36070 7200 36100 7440
rect 28700 7170 36100 7200
rect 28700 6930 28780 7170
rect 29020 6930 29110 7170
rect 29350 6930 29440 7170
rect 29680 6930 29770 7170
rect 30010 6930 30100 7170
rect 30340 6930 30430 7170
rect 30670 6930 30760 7170
rect 31000 6930 31090 7170
rect 31330 6930 31420 7170
rect 31660 6930 31750 7170
rect 31990 6930 32080 7170
rect 32320 6930 32410 7170
rect 32650 6930 32740 7170
rect 32980 6930 33070 7170
rect 33310 6930 33400 7170
rect 33640 6930 33730 7170
rect 33970 6930 34060 7170
rect 34300 6930 34390 7170
rect 34630 6930 34720 7170
rect 34960 6930 35050 7170
rect 35290 7070 36100 7170
rect 35290 6930 35830 7070
rect 28700 6840 35830 6930
rect 28700 6600 28780 6840
rect 29020 6600 29110 6840
rect 29350 6600 29440 6840
rect 29680 6600 29770 6840
rect 30010 6600 30100 6840
rect 30340 6600 30430 6840
rect 30670 6600 30760 6840
rect 31000 6600 31090 6840
rect 31330 6600 31420 6840
rect 31660 6600 31750 6840
rect 31990 6600 32080 6840
rect 32320 6600 32410 6840
rect 32650 6600 32740 6840
rect 32980 6600 33070 6840
rect 33310 6600 33400 6840
rect 33640 6600 33730 6840
rect 33970 6600 34060 6840
rect 34300 6600 34390 6840
rect 34630 6600 34720 6840
rect 34960 6600 35050 6840
rect 35290 6830 35830 6840
rect 36070 6830 36100 7070
rect 35290 6740 36100 6830
rect 35290 6600 35830 6740
rect 28700 6510 35830 6600
rect 28700 6270 28780 6510
rect 29020 6270 29110 6510
rect 29350 6270 29440 6510
rect 29680 6270 29770 6510
rect 30010 6270 30100 6510
rect 30340 6270 30430 6510
rect 30670 6270 30760 6510
rect 31000 6270 31090 6510
rect 31330 6270 31420 6510
rect 31660 6270 31750 6510
rect 31990 6270 32080 6510
rect 32320 6270 32410 6510
rect 32650 6270 32740 6510
rect 32980 6270 33070 6510
rect 33310 6270 33400 6510
rect 33640 6270 33730 6510
rect 33970 6270 34060 6510
rect 34300 6270 34390 6510
rect 34630 6270 34720 6510
rect 34960 6270 35050 6510
rect 35290 6500 35830 6510
rect 36070 6500 36100 6740
rect 35290 6410 36100 6500
rect 35290 6270 35830 6410
rect 28700 6180 35830 6270
rect 28700 5940 28780 6180
rect 29020 5940 29110 6180
rect 29350 5940 29440 6180
rect 29680 5940 29770 6180
rect 30010 5940 30100 6180
rect 30340 5940 30430 6180
rect 30670 5940 30760 6180
rect 31000 5940 31090 6180
rect 31330 5940 31420 6180
rect 31660 5940 31750 6180
rect 31990 5940 32080 6180
rect 32320 5940 32410 6180
rect 32650 5940 32740 6180
rect 32980 5940 33070 6180
rect 33310 5940 33400 6180
rect 33640 5940 33730 6180
rect 33970 5940 34060 6180
rect 34300 5940 34390 6180
rect 34630 5940 34720 6180
rect 34960 5940 35050 6180
rect 35290 6170 35830 6180
rect 36070 6170 36100 6410
rect 35290 6080 36100 6170
rect 35290 5940 35830 6080
rect 28700 5850 35830 5940
rect 28700 5610 28780 5850
rect 29020 5610 29110 5850
rect 29350 5610 29440 5850
rect 29680 5610 29770 5850
rect 30010 5610 30100 5850
rect 30340 5610 30430 5850
rect 30670 5610 30760 5850
rect 31000 5610 31090 5850
rect 31330 5610 31420 5850
rect 31660 5610 31750 5850
rect 31990 5610 32080 5850
rect 32320 5610 32410 5850
rect 32650 5610 32740 5850
rect 32980 5610 33070 5850
rect 33310 5610 33400 5850
rect 33640 5610 33730 5850
rect 33970 5610 34060 5850
rect 34300 5610 34390 5850
rect 34630 5610 34720 5850
rect 34960 5610 35050 5850
rect 35290 5840 35830 5850
rect 36070 5840 36100 6080
rect 35290 5750 36100 5840
rect 35290 5610 35830 5750
rect 28700 5520 35830 5610
rect 28700 5280 28780 5520
rect 29020 5280 29110 5520
rect 29350 5280 29440 5520
rect 29680 5280 29770 5520
rect 30010 5280 30100 5520
rect 30340 5280 30430 5520
rect 30670 5280 30760 5520
rect 31000 5280 31090 5520
rect 31330 5280 31420 5520
rect 31660 5280 31750 5520
rect 31990 5280 32080 5520
rect 32320 5280 32410 5520
rect 32650 5280 32740 5520
rect 32980 5280 33070 5520
rect 33310 5280 33400 5520
rect 33640 5280 33730 5520
rect 33970 5280 34060 5520
rect 34300 5280 34390 5520
rect 34630 5280 34720 5520
rect 34960 5280 35050 5520
rect 35290 5510 35830 5520
rect 36070 5510 36100 5750
rect 35290 5420 36100 5510
rect 35290 5280 35830 5420
rect 28700 5190 35830 5280
rect 28700 4950 28780 5190
rect 29020 4950 29110 5190
rect 29350 4950 29440 5190
rect 29680 4950 29770 5190
rect 30010 4950 30100 5190
rect 30340 4950 30430 5190
rect 30670 4950 30760 5190
rect 31000 4950 31090 5190
rect 31330 4950 31420 5190
rect 31660 4950 31750 5190
rect 31990 4950 32080 5190
rect 32320 4950 32410 5190
rect 32650 4950 32740 5190
rect 32980 4950 33070 5190
rect 33310 4950 33400 5190
rect 33640 4950 33730 5190
rect 33970 4950 34060 5190
rect 34300 4950 34390 5190
rect 34630 4950 34720 5190
rect 34960 4950 35050 5190
rect 35290 5180 35830 5190
rect 36070 5180 36100 5420
rect 35290 5090 36100 5180
rect 35290 4950 35830 5090
rect 28700 4860 35830 4950
rect 28700 4620 28780 4860
rect 29020 4620 29110 4860
rect 29350 4620 29440 4860
rect 29680 4620 29770 4860
rect 30010 4620 30100 4860
rect 30340 4620 30430 4860
rect 30670 4620 30760 4860
rect 31000 4620 31090 4860
rect 31330 4620 31420 4860
rect 31660 4620 31750 4860
rect 31990 4620 32080 4860
rect 32320 4620 32410 4860
rect 32650 4620 32740 4860
rect 32980 4620 33070 4860
rect 33310 4620 33400 4860
rect 33640 4620 33730 4860
rect 33970 4620 34060 4860
rect 34300 4620 34390 4860
rect 34630 4620 34720 4860
rect 34960 4620 35050 4860
rect 35290 4850 35830 4860
rect 36070 4850 36100 5090
rect 35290 4760 36100 4850
rect 35290 4620 35830 4760
rect 28700 4530 35830 4620
rect 28700 4290 28780 4530
rect 29020 4290 29110 4530
rect 29350 4290 29440 4530
rect 29680 4290 29770 4530
rect 30010 4290 30100 4530
rect 30340 4290 30430 4530
rect 30670 4290 30760 4530
rect 31000 4290 31090 4530
rect 31330 4290 31420 4530
rect 31660 4290 31750 4530
rect 31990 4290 32080 4530
rect 32320 4290 32410 4530
rect 32650 4290 32740 4530
rect 32980 4290 33070 4530
rect 33310 4290 33400 4530
rect 33640 4290 33730 4530
rect 33970 4290 34060 4530
rect 34300 4290 34390 4530
rect 34630 4290 34720 4530
rect 34960 4290 35050 4530
rect 35290 4520 35830 4530
rect 36070 4520 36100 4760
rect 35290 4430 36100 4520
rect 35290 4290 35830 4430
rect 28700 4200 35830 4290
rect 28700 3960 28780 4200
rect 29020 3960 29110 4200
rect 29350 3960 29440 4200
rect 29680 3960 29770 4200
rect 30010 3960 30100 4200
rect 30340 3960 30430 4200
rect 30670 3960 30760 4200
rect 31000 3960 31090 4200
rect 31330 3960 31420 4200
rect 31660 3960 31750 4200
rect 31990 3960 32080 4200
rect 32320 3960 32410 4200
rect 32650 3960 32740 4200
rect 32980 3960 33070 4200
rect 33310 3960 33400 4200
rect 33640 3960 33730 4200
rect 33970 3960 34060 4200
rect 34300 3960 34390 4200
rect 34630 3960 34720 4200
rect 34960 3960 35050 4200
rect 35290 4190 35830 4200
rect 36070 4190 36100 4430
rect 35290 4060 36100 4190
rect 35290 3960 35830 4060
rect 28700 3870 35830 3960
rect 28700 3630 28780 3870
rect 29020 3630 29110 3870
rect 29350 3630 29440 3870
rect 29680 3630 29770 3870
rect 30010 3630 30100 3870
rect 30340 3630 30430 3870
rect 30670 3630 30760 3870
rect 31000 3630 31090 3870
rect 31330 3630 31420 3870
rect 31660 3630 31750 3870
rect 31990 3630 32080 3870
rect 32320 3630 32410 3870
rect 32650 3630 32740 3870
rect 32980 3630 33070 3870
rect 33310 3630 33400 3870
rect 33640 3630 33730 3870
rect 33970 3630 34060 3870
rect 34300 3630 34390 3870
rect 34630 3630 34720 3870
rect 34960 3630 35050 3870
rect 35290 3820 35830 3870
rect 36070 3820 36100 4060
rect 35290 3730 36100 3820
rect 35290 3630 35830 3730
rect 28700 3540 35830 3630
rect 28700 3300 28780 3540
rect 29020 3300 29110 3540
rect 29350 3300 29440 3540
rect 29680 3300 29770 3540
rect 30010 3300 30100 3540
rect 30340 3300 30430 3540
rect 30670 3300 30760 3540
rect 31000 3300 31090 3540
rect 31330 3300 31420 3540
rect 31660 3300 31750 3540
rect 31990 3300 32080 3540
rect 32320 3300 32410 3540
rect 32650 3300 32740 3540
rect 32980 3300 33070 3540
rect 33310 3300 33400 3540
rect 33640 3300 33730 3540
rect 33970 3300 34060 3540
rect 34300 3300 34390 3540
rect 34630 3300 34720 3540
rect 34960 3300 35050 3540
rect 35290 3490 35830 3540
rect 36070 3490 36100 3730
rect 35290 3400 36100 3490
rect 35290 3300 35830 3400
rect 28700 3210 35830 3300
rect 28700 2970 28780 3210
rect 29020 2970 29110 3210
rect 29350 2970 29440 3210
rect 29680 2970 29770 3210
rect 30010 2970 30100 3210
rect 30340 2970 30430 3210
rect 30670 2970 30760 3210
rect 31000 2970 31090 3210
rect 31330 2970 31420 3210
rect 31660 2970 31750 3210
rect 31990 2970 32080 3210
rect 32320 2970 32410 3210
rect 32650 2970 32740 3210
rect 32980 2970 33070 3210
rect 33310 2970 33400 3210
rect 33640 2970 33730 3210
rect 33970 2970 34060 3210
rect 34300 2970 34390 3210
rect 34630 2970 34720 3210
rect 34960 2970 35050 3210
rect 35290 3160 35830 3210
rect 36070 3160 36100 3400
rect 35290 3070 36100 3160
rect 35290 2970 35830 3070
rect 28700 2880 35830 2970
rect 28700 2640 28780 2880
rect 29020 2640 29110 2880
rect 29350 2640 29440 2880
rect 29680 2640 29770 2880
rect 30010 2640 30100 2880
rect 30340 2640 30430 2880
rect 30670 2640 30760 2880
rect 31000 2640 31090 2880
rect 31330 2640 31420 2880
rect 31660 2640 31750 2880
rect 31990 2640 32080 2880
rect 32320 2640 32410 2880
rect 32650 2640 32740 2880
rect 32980 2640 33070 2880
rect 33310 2640 33400 2880
rect 33640 2640 33730 2880
rect 33970 2640 34060 2880
rect 34300 2640 34390 2880
rect 34630 2640 34720 2880
rect 34960 2640 35050 2880
rect 35290 2830 35830 2880
rect 36070 2830 36100 3070
rect 35290 2740 36100 2830
rect 35290 2640 35830 2740
rect 28700 2550 35830 2640
rect 28700 2310 28780 2550
rect 29020 2310 29110 2550
rect 29350 2310 29440 2550
rect 29680 2310 29770 2550
rect 30010 2310 30100 2550
rect 30340 2310 30430 2550
rect 30670 2310 30760 2550
rect 31000 2310 31090 2550
rect 31330 2310 31420 2550
rect 31660 2310 31750 2550
rect 31990 2310 32080 2550
rect 32320 2310 32410 2550
rect 32650 2310 32740 2550
rect 32980 2310 33070 2550
rect 33310 2310 33400 2550
rect 33640 2310 33730 2550
rect 33970 2310 34060 2550
rect 34300 2310 34390 2550
rect 34630 2310 34720 2550
rect 34960 2310 35050 2550
rect 35290 2500 35830 2550
rect 36070 2500 36100 2740
rect 35290 2410 36100 2500
rect 35290 2310 35830 2410
rect 28700 2220 35830 2310
rect 28700 1980 28780 2220
rect 29020 1980 29110 2220
rect 29350 1980 29440 2220
rect 29680 1980 29770 2220
rect 30010 1980 30100 2220
rect 30340 1980 30430 2220
rect 30670 1980 30760 2220
rect 31000 1980 31090 2220
rect 31330 1980 31420 2220
rect 31660 1980 31750 2220
rect 31990 1980 32080 2220
rect 32320 1980 32410 2220
rect 32650 1980 32740 2220
rect 32980 1980 33070 2220
rect 33310 1980 33400 2220
rect 33640 1980 33730 2220
rect 33970 1980 34060 2220
rect 34300 1980 34390 2220
rect 34630 1980 34720 2220
rect 34960 1980 35050 2220
rect 35290 2170 35830 2220
rect 36070 2170 36100 2410
rect 35290 2080 36100 2170
rect 35290 1980 35830 2080
rect 28700 1890 35830 1980
rect 28700 1650 28780 1890
rect 29020 1650 29110 1890
rect 29350 1650 29440 1890
rect 29680 1650 29770 1890
rect 30010 1650 30100 1890
rect 30340 1650 30430 1890
rect 30670 1650 30760 1890
rect 31000 1650 31090 1890
rect 31330 1650 31420 1890
rect 31660 1650 31750 1890
rect 31990 1650 32080 1890
rect 32320 1650 32410 1890
rect 32650 1650 32740 1890
rect 32980 1650 33070 1890
rect 33310 1650 33400 1890
rect 33640 1650 33730 1890
rect 33970 1650 34060 1890
rect 34300 1650 34390 1890
rect 34630 1650 34720 1890
rect 34960 1650 35050 1890
rect 35290 1840 35830 1890
rect 36070 1840 36100 2080
rect 35290 1750 36100 1840
rect 35290 1650 35830 1750
rect 28700 1560 35830 1650
rect 28700 1320 28780 1560
rect 29020 1320 29110 1560
rect 29350 1320 29440 1560
rect 29680 1320 29770 1560
rect 30010 1320 30100 1560
rect 30340 1320 30430 1560
rect 30670 1320 30760 1560
rect 31000 1320 31090 1560
rect 31330 1320 31420 1560
rect 31660 1320 31750 1560
rect 31990 1320 32080 1560
rect 32320 1320 32410 1560
rect 32650 1320 32740 1560
rect 32980 1320 33070 1560
rect 33310 1320 33400 1560
rect 33640 1320 33730 1560
rect 33970 1320 34060 1560
rect 34300 1320 34390 1560
rect 34630 1320 34720 1560
rect 34960 1320 35050 1560
rect 35290 1510 35830 1560
rect 36070 1510 36100 1750
rect 35290 1420 36100 1510
rect 35290 1320 35830 1420
rect 28700 1180 35830 1320
rect 36070 1180 36100 1420
rect 21060 980 21540 1040
rect 21060 740 21110 980
rect 21480 740 21540 980
rect 21060 710 21540 740
rect 23460 980 23940 1040
rect 23460 740 23510 980
rect 23880 740 23940 980
rect 23460 710 23940 740
rect -170 -1840 19210 -1040
rect -6530 -2720 14530 -2160
rect -6530 -2960 1720 -2720
rect 1960 -2960 2050 -2720
rect 2290 -2960 2390 -2720
rect 2630 -2960 2720 -2720
rect 2960 -2960 11940 -2720
rect 12180 -2960 12270 -2720
rect 12510 -2960 12610 -2720
rect 12850 -2960 12940 -2720
rect 13180 -2960 14530 -2720
rect -6530 -11680 -2530 -2960
rect 1540 -2990 3140 -2960
rect 11760 -2990 13360 -2960
rect 15210 -3840 19210 -1840
rect 28700 230 36100 1180
rect 28700 -10 28780 230
rect 29020 -10 29110 230
rect 29350 -10 29440 230
rect 29680 -10 29770 230
rect 30010 -10 30100 230
rect 30340 -10 30430 230
rect 30670 -10 30760 230
rect 31000 -10 31090 230
rect 31330 -10 31420 230
rect 31660 -10 31750 230
rect 31990 -10 32080 230
rect 32320 -10 32410 230
rect 32650 -10 32740 230
rect 32980 -10 33070 230
rect 33310 -10 33400 230
rect 33640 -10 33730 230
rect 33970 -10 34060 230
rect 34300 -10 34390 230
rect 34630 -10 34720 230
rect 34960 -10 35050 230
rect 35290 170 36100 230
rect 35290 -10 35830 170
rect 28700 -70 35830 -10
rect 36070 -70 36100 170
rect 28700 -100 36100 -70
rect 28700 -340 28780 -100
rect 29020 -340 29110 -100
rect 29350 -340 29440 -100
rect 29680 -340 29770 -100
rect 30010 -340 30100 -100
rect 30340 -340 30430 -100
rect 30670 -340 30760 -100
rect 31000 -340 31090 -100
rect 31330 -340 31420 -100
rect 31660 -340 31750 -100
rect 31990 -340 32080 -100
rect 32320 -340 32410 -100
rect 32650 -340 32740 -100
rect 32980 -340 33070 -100
rect 33310 -340 33400 -100
rect 33640 -340 33730 -100
rect 33970 -340 34060 -100
rect 34300 -340 34390 -100
rect 34630 -340 34720 -100
rect 34960 -340 35050 -100
rect 35290 -160 36100 -100
rect 35290 -340 35830 -160
rect 28700 -400 35830 -340
rect 36070 -400 36100 -160
rect 28700 -430 36100 -400
rect 28700 -670 28780 -430
rect 29020 -670 29110 -430
rect 29350 -670 29440 -430
rect 29680 -670 29770 -430
rect 30010 -670 30100 -430
rect 30340 -670 30430 -430
rect 30670 -670 30760 -430
rect 31000 -670 31090 -430
rect 31330 -670 31420 -430
rect 31660 -670 31750 -430
rect 31990 -670 32080 -430
rect 32320 -670 32410 -430
rect 32650 -670 32740 -430
rect 32980 -670 33070 -430
rect 33310 -670 33400 -430
rect 33640 -670 33730 -430
rect 33970 -670 34060 -430
rect 34300 -670 34390 -430
rect 34630 -670 34720 -430
rect 34960 -670 35050 -430
rect 35290 -530 36100 -430
rect 35290 -670 35830 -530
rect 28700 -760 35830 -670
rect 28700 -1000 28780 -760
rect 29020 -1000 29110 -760
rect 29350 -1000 29440 -760
rect 29680 -1000 29770 -760
rect 30010 -1000 30100 -760
rect 30340 -1000 30430 -760
rect 30670 -1000 30760 -760
rect 31000 -1000 31090 -760
rect 31330 -1000 31420 -760
rect 31660 -1000 31750 -760
rect 31990 -1000 32080 -760
rect 32320 -1000 32410 -760
rect 32650 -1000 32740 -760
rect 32980 -1000 33070 -760
rect 33310 -1000 33400 -760
rect 33640 -1000 33730 -760
rect 33970 -1000 34060 -760
rect 34300 -1000 34390 -760
rect 34630 -1000 34720 -760
rect 34960 -1000 35050 -760
rect 35290 -770 35830 -760
rect 36070 -770 36100 -530
rect 35290 -860 36100 -770
rect 35290 -1000 35830 -860
rect 28700 -1090 35830 -1000
rect 28700 -1330 28780 -1090
rect 29020 -1330 29110 -1090
rect 29350 -1330 29440 -1090
rect 29680 -1330 29770 -1090
rect 30010 -1330 30100 -1090
rect 30340 -1330 30430 -1090
rect 30670 -1330 30760 -1090
rect 31000 -1330 31090 -1090
rect 31330 -1330 31420 -1090
rect 31660 -1330 31750 -1090
rect 31990 -1330 32080 -1090
rect 32320 -1330 32410 -1090
rect 32650 -1330 32740 -1090
rect 32980 -1330 33070 -1090
rect 33310 -1330 33400 -1090
rect 33640 -1330 33730 -1090
rect 33970 -1330 34060 -1090
rect 34300 -1330 34390 -1090
rect 34630 -1330 34720 -1090
rect 34960 -1330 35050 -1090
rect 35290 -1100 35830 -1090
rect 36070 -1100 36100 -860
rect 35290 -1190 36100 -1100
rect 35290 -1330 35830 -1190
rect 28700 -1420 35830 -1330
rect 28700 -1660 28780 -1420
rect 29020 -1660 29110 -1420
rect 29350 -1660 29440 -1420
rect 29680 -1660 29770 -1420
rect 30010 -1660 30100 -1420
rect 30340 -1660 30430 -1420
rect 30670 -1660 30760 -1420
rect 31000 -1660 31090 -1420
rect 31330 -1660 31420 -1420
rect 31660 -1660 31750 -1420
rect 31990 -1660 32080 -1420
rect 32320 -1660 32410 -1420
rect 32650 -1660 32740 -1420
rect 32980 -1660 33070 -1420
rect 33310 -1660 33400 -1420
rect 33640 -1660 33730 -1420
rect 33970 -1660 34060 -1420
rect 34300 -1660 34390 -1420
rect 34630 -1660 34720 -1420
rect 34960 -1660 35050 -1420
rect 35290 -1430 35830 -1420
rect 36070 -1430 36100 -1190
rect 35290 -1520 36100 -1430
rect 35290 -1660 35830 -1520
rect 28700 -1750 35830 -1660
rect 28700 -1990 28780 -1750
rect 29020 -1990 29110 -1750
rect 29350 -1990 29440 -1750
rect 29680 -1990 29770 -1750
rect 30010 -1990 30100 -1750
rect 30340 -1990 30430 -1750
rect 30670 -1990 30760 -1750
rect 31000 -1990 31090 -1750
rect 31330 -1990 31420 -1750
rect 31660 -1990 31750 -1750
rect 31990 -1990 32080 -1750
rect 32320 -1990 32410 -1750
rect 32650 -1990 32740 -1750
rect 32980 -1990 33070 -1750
rect 33310 -1990 33400 -1750
rect 33640 -1990 33730 -1750
rect 33970 -1990 34060 -1750
rect 34300 -1990 34390 -1750
rect 34630 -1990 34720 -1750
rect 34960 -1990 35050 -1750
rect 35290 -1760 35830 -1750
rect 36070 -1760 36100 -1520
rect 35290 -1850 36100 -1760
rect 35290 -1990 35830 -1850
rect 28700 -2080 35830 -1990
rect 28700 -2320 28780 -2080
rect 29020 -2320 29110 -2080
rect 29350 -2320 29440 -2080
rect 29680 -2320 29770 -2080
rect 30010 -2320 30100 -2080
rect 30340 -2320 30430 -2080
rect 30670 -2320 30760 -2080
rect 31000 -2320 31090 -2080
rect 31330 -2320 31420 -2080
rect 31660 -2320 31750 -2080
rect 31990 -2320 32080 -2080
rect 32320 -2320 32410 -2080
rect 32650 -2320 32740 -2080
rect 32980 -2320 33070 -2080
rect 33310 -2320 33400 -2080
rect 33640 -2320 33730 -2080
rect 33970 -2320 34060 -2080
rect 34300 -2320 34390 -2080
rect 34630 -2320 34720 -2080
rect 34960 -2320 35050 -2080
rect 35290 -2090 35830 -2080
rect 36070 -2090 36100 -1850
rect 35290 -2180 36100 -2090
rect 35290 -2320 35830 -2180
rect 28700 -2410 35830 -2320
rect 28700 -2650 28780 -2410
rect 29020 -2650 29110 -2410
rect 29350 -2650 29440 -2410
rect 29680 -2650 29770 -2410
rect 30010 -2650 30100 -2410
rect 30340 -2650 30430 -2410
rect 30670 -2650 30760 -2410
rect 31000 -2650 31090 -2410
rect 31330 -2650 31420 -2410
rect 31660 -2650 31750 -2410
rect 31990 -2650 32080 -2410
rect 32320 -2650 32410 -2410
rect 32650 -2650 32740 -2410
rect 32980 -2650 33070 -2410
rect 33310 -2650 33400 -2410
rect 33640 -2650 33730 -2410
rect 33970 -2650 34060 -2410
rect 34300 -2650 34390 -2410
rect 34630 -2650 34720 -2410
rect 34960 -2650 35050 -2410
rect 35290 -2420 35830 -2410
rect 36070 -2420 36100 -2180
rect 35290 -2510 36100 -2420
rect 35290 -2650 35830 -2510
rect 28700 -2740 35830 -2650
rect 28700 -2980 28780 -2740
rect 29020 -2980 29110 -2740
rect 29350 -2980 29440 -2740
rect 29680 -2980 29770 -2740
rect 30010 -2980 30100 -2740
rect 30340 -2980 30430 -2740
rect 30670 -2980 30760 -2740
rect 31000 -2980 31090 -2740
rect 31330 -2980 31420 -2740
rect 31660 -2980 31750 -2740
rect 31990 -2980 32080 -2740
rect 32320 -2980 32410 -2740
rect 32650 -2980 32740 -2740
rect 32980 -2980 33070 -2740
rect 33310 -2980 33400 -2740
rect 33640 -2980 33730 -2740
rect 33970 -2980 34060 -2740
rect 34300 -2980 34390 -2740
rect 34630 -2980 34720 -2740
rect 34960 -2980 35050 -2740
rect 35290 -2750 35830 -2740
rect 36070 -2750 36100 -2510
rect 35290 -2840 36100 -2750
rect 35290 -2980 35830 -2840
rect 28700 -3070 35830 -2980
rect 28700 -3310 28780 -3070
rect 29020 -3310 29110 -3070
rect 29350 -3310 29440 -3070
rect 29680 -3310 29770 -3070
rect 30010 -3310 30100 -3070
rect 30340 -3310 30430 -3070
rect 30670 -3310 30760 -3070
rect 31000 -3310 31090 -3070
rect 31330 -3310 31420 -3070
rect 31660 -3310 31750 -3070
rect 31990 -3310 32080 -3070
rect 32320 -3310 32410 -3070
rect 32650 -3310 32740 -3070
rect 32980 -3310 33070 -3070
rect 33310 -3310 33400 -3070
rect 33640 -3310 33730 -3070
rect 33970 -3310 34060 -3070
rect 34300 -3310 34390 -3070
rect 34630 -3310 34720 -3070
rect 34960 -3310 35050 -3070
rect 35290 -3080 35830 -3070
rect 36070 -3080 36100 -2840
rect 35290 -3170 36100 -3080
rect 35290 -3310 35830 -3170
rect 28700 -3400 35830 -3310
rect 28700 -3640 28780 -3400
rect 29020 -3640 29110 -3400
rect 29350 -3640 29440 -3400
rect 29680 -3640 29770 -3400
rect 30010 -3640 30100 -3400
rect 30340 -3640 30430 -3400
rect 30670 -3640 30760 -3400
rect 31000 -3640 31090 -3400
rect 31330 -3640 31420 -3400
rect 31660 -3640 31750 -3400
rect 31990 -3640 32080 -3400
rect 32320 -3640 32410 -3400
rect 32650 -3640 32740 -3400
rect 32980 -3640 33070 -3400
rect 33310 -3640 33400 -3400
rect 33640 -3640 33730 -3400
rect 33970 -3640 34060 -3400
rect 34300 -3640 34390 -3400
rect 34630 -3640 34720 -3400
rect 34960 -3640 35050 -3400
rect 35290 -3410 35830 -3400
rect 36070 -3410 36100 -3170
rect 35290 -3540 36100 -3410
rect 35290 -3640 35830 -3540
rect 20020 -3690 20500 -3660
rect 20020 -3840 20080 -3690
rect 15210 -3930 20080 -3840
rect 20450 -3840 20500 -3690
rect 24500 -3690 24980 -3660
rect 24500 -3840 24560 -3690
rect 20450 -3930 24560 -3840
rect 24930 -3840 24980 -3690
rect 28700 -3730 35830 -3640
rect 28700 -3840 28780 -3730
rect 24930 -3850 26820 -3840
rect 27980 -3850 28780 -3840
rect 24930 -3930 28780 -3850
rect 15210 -3970 28780 -3930
rect 29020 -3970 29110 -3730
rect 29350 -3970 29440 -3730
rect 29680 -3970 29770 -3730
rect 30010 -3970 30100 -3730
rect 30340 -3970 30430 -3730
rect 30670 -3970 30760 -3730
rect 31000 -3970 31090 -3730
rect 31330 -3970 31420 -3730
rect 31660 -3970 31750 -3730
rect 31990 -3970 32080 -3730
rect 32320 -3970 32410 -3730
rect 32650 -3970 32740 -3730
rect 32980 -3970 33070 -3730
rect 33310 -3970 33400 -3730
rect 33640 -3970 33730 -3730
rect 33970 -3970 34060 -3730
rect 34300 -3970 34390 -3730
rect 34630 -3970 34720 -3730
rect 34960 -3970 35050 -3730
rect 35290 -3780 35830 -3730
rect 36070 -3780 36100 -3540
rect 35290 -3870 36100 -3780
rect 35290 -3970 35830 -3870
rect -1860 -4250 150 -4050
rect -1860 -4260 -120 -4250
rect -1860 -4500 -1650 -4260
rect -1410 -4500 -1320 -4260
rect -1080 -4500 -990 -4260
rect -750 -4500 -660 -4260
rect -420 -4490 -120 -4260
rect 120 -4490 150 -4250
rect -420 -4500 150 -4490
rect -1860 -4580 150 -4500
rect -1860 -4590 -120 -4580
rect -1860 -4830 -1650 -4590
rect -1410 -4830 -1320 -4590
rect -1080 -4830 -990 -4590
rect -750 -4830 -660 -4590
rect -420 -4820 -120 -4590
rect 120 -4820 150 -4580
rect -420 -4830 150 -4820
rect -1860 -4910 150 -4830
rect -1860 -4920 -120 -4910
rect -1860 -5160 -1650 -4920
rect -1410 -5160 -1320 -4920
rect -1080 -5160 -990 -4920
rect -750 -5160 -660 -4920
rect -420 -5150 -120 -4920
rect 120 -5150 150 -4910
rect -420 -5160 150 -5150
rect -1860 -5240 150 -5160
rect -1860 -5250 -120 -5240
rect -1860 -5490 -1650 -5250
rect -1410 -5490 -1320 -5250
rect -1080 -5490 -990 -5250
rect -750 -5490 -660 -5250
rect -420 -5480 -120 -5250
rect 120 -5480 150 -5240
rect -420 -5490 150 -5480
rect -1860 -5660 150 -5490
rect 15210 -4060 35830 -3970
rect 15210 -4240 28780 -4060
rect -1860 -7650 150 -7450
rect -1860 -7660 -120 -7650
rect -1860 -7900 -1650 -7660
rect -1410 -7900 -1320 -7660
rect -1080 -7900 -990 -7660
rect -750 -7900 -660 -7660
rect -420 -7890 -120 -7660
rect 120 -7890 150 -7650
rect -420 -7900 150 -7890
rect -1860 -7980 150 -7900
rect -1860 -7990 -120 -7980
rect -1860 -8230 -1650 -7990
rect -1410 -8230 -1320 -7990
rect -1080 -8230 -990 -7990
rect -750 -8230 -660 -7990
rect -420 -8220 -120 -7990
rect 120 -8220 150 -7980
rect -420 -8230 150 -8220
rect -1860 -8310 150 -8230
rect -1860 -8320 -120 -8310
rect -1860 -8560 -1650 -8320
rect -1410 -8560 -1320 -8320
rect -1080 -8560 -990 -8320
rect -750 -8560 -660 -8320
rect -420 -8550 -120 -8320
rect 120 -8550 150 -8310
rect -420 -8560 150 -8550
rect -1860 -8640 150 -8560
rect -1860 -8650 -120 -8640
rect -1860 -8890 -1650 -8650
rect -1410 -8890 -1320 -8650
rect -1080 -8890 -990 -8650
rect -750 -8890 -660 -8650
rect -420 -8880 -120 -8650
rect 120 -8880 150 -8640
rect -420 -8890 150 -8880
rect -1860 -9060 150 -8890
rect 15210 -8530 19210 -4240
rect 26820 -4250 27980 -4240
rect 28700 -4300 28780 -4240
rect 29020 -4300 29110 -4060
rect 29350 -4300 29440 -4060
rect 29680 -4300 29770 -4060
rect 30010 -4300 30100 -4060
rect 30340 -4300 30430 -4060
rect 30670 -4300 30760 -4060
rect 31000 -4300 31090 -4060
rect 31330 -4300 31420 -4060
rect 31660 -4300 31750 -4060
rect 31990 -4300 32080 -4060
rect 32320 -4300 32410 -4060
rect 32650 -4300 32740 -4060
rect 32980 -4300 33070 -4060
rect 33310 -4300 33400 -4060
rect 33640 -4300 33730 -4060
rect 33970 -4300 34060 -4060
rect 34300 -4300 34390 -4060
rect 34630 -4300 34720 -4060
rect 34960 -4300 35050 -4060
rect 35290 -4110 35830 -4060
rect 36070 -4110 36100 -3870
rect 35290 -4200 36100 -4110
rect 35290 -4300 35830 -4200
rect 28700 -4390 35830 -4300
rect 28700 -4630 28780 -4390
rect 29020 -4630 29110 -4390
rect 29350 -4630 29440 -4390
rect 29680 -4630 29770 -4390
rect 30010 -4630 30100 -4390
rect 30340 -4630 30430 -4390
rect 30670 -4630 30760 -4390
rect 31000 -4630 31090 -4390
rect 31330 -4630 31420 -4390
rect 31660 -4630 31750 -4390
rect 31990 -4630 32080 -4390
rect 32320 -4630 32410 -4390
rect 32650 -4630 32740 -4390
rect 32980 -4630 33070 -4390
rect 33310 -4630 33400 -4390
rect 33640 -4630 33730 -4390
rect 33970 -4630 34060 -4390
rect 34300 -4630 34390 -4390
rect 34630 -4630 34720 -4390
rect 34960 -4630 35050 -4390
rect 35290 -4440 35830 -4390
rect 36070 -4440 36100 -4200
rect 35290 -4530 36100 -4440
rect 35290 -4630 35830 -4530
rect 28700 -4720 35830 -4630
rect 28700 -4960 28780 -4720
rect 29020 -4960 29110 -4720
rect 29350 -4960 29440 -4720
rect 29680 -4960 29770 -4720
rect 30010 -4960 30100 -4720
rect 30340 -4960 30430 -4720
rect 30670 -4960 30760 -4720
rect 31000 -4960 31090 -4720
rect 31330 -4960 31420 -4720
rect 31660 -4960 31750 -4720
rect 31990 -4960 32080 -4720
rect 32320 -4960 32410 -4720
rect 32650 -4960 32740 -4720
rect 32980 -4960 33070 -4720
rect 33310 -4960 33400 -4720
rect 33640 -4960 33730 -4720
rect 33970 -4960 34060 -4720
rect 34300 -4960 34390 -4720
rect 34630 -4960 34720 -4720
rect 34960 -4960 35050 -4720
rect 35290 -4770 35830 -4720
rect 36070 -4770 36100 -4530
rect 35290 -4860 36100 -4770
rect 35290 -4960 35830 -4860
rect 28700 -5050 35830 -4960
rect 28700 -5290 28780 -5050
rect 29020 -5290 29110 -5050
rect 29350 -5290 29440 -5050
rect 29680 -5290 29770 -5050
rect 30010 -5290 30100 -5050
rect 30340 -5290 30430 -5050
rect 30670 -5290 30760 -5050
rect 31000 -5290 31090 -5050
rect 31330 -5290 31420 -5050
rect 31660 -5290 31750 -5050
rect 31990 -5290 32080 -5050
rect 32320 -5290 32410 -5050
rect 32650 -5290 32740 -5050
rect 32980 -5290 33070 -5050
rect 33310 -5290 33400 -5050
rect 33640 -5290 33730 -5050
rect 33970 -5290 34060 -5050
rect 34300 -5290 34390 -5050
rect 34630 -5290 34720 -5050
rect 34960 -5290 35050 -5050
rect 35290 -5100 35830 -5050
rect 36070 -5100 36100 -4860
rect 35290 -5190 36100 -5100
rect 35290 -5290 35830 -5190
rect 28700 -5380 35830 -5290
rect 28700 -5620 28780 -5380
rect 29020 -5620 29110 -5380
rect 29350 -5620 29440 -5380
rect 29680 -5620 29770 -5380
rect 30010 -5620 30100 -5380
rect 30340 -5620 30430 -5380
rect 30670 -5620 30760 -5380
rect 31000 -5620 31090 -5380
rect 31330 -5620 31420 -5380
rect 31660 -5620 31750 -5380
rect 31990 -5620 32080 -5380
rect 32320 -5620 32410 -5380
rect 32650 -5620 32740 -5380
rect 32980 -5620 33070 -5380
rect 33310 -5620 33400 -5380
rect 33640 -5620 33730 -5380
rect 33970 -5620 34060 -5380
rect 34300 -5620 34390 -5380
rect 34630 -5620 34720 -5380
rect 34960 -5620 35050 -5380
rect 35290 -5430 35830 -5380
rect 36070 -5430 36100 -5190
rect 35290 -5520 36100 -5430
rect 35290 -5620 35830 -5520
rect 28700 -5710 35830 -5620
rect 28700 -5950 28780 -5710
rect 29020 -5950 29110 -5710
rect 29350 -5950 29440 -5710
rect 29680 -5950 29770 -5710
rect 30010 -5950 30100 -5710
rect 30340 -5950 30430 -5710
rect 30670 -5950 30760 -5710
rect 31000 -5950 31090 -5710
rect 31330 -5950 31420 -5710
rect 31660 -5950 31750 -5710
rect 31990 -5950 32080 -5710
rect 32320 -5950 32410 -5710
rect 32650 -5950 32740 -5710
rect 32980 -5950 33070 -5710
rect 33310 -5950 33400 -5710
rect 33640 -5950 33730 -5710
rect 33970 -5950 34060 -5710
rect 34300 -5950 34390 -5710
rect 34630 -5950 34720 -5710
rect 34960 -5950 35050 -5710
rect 35290 -5760 35830 -5710
rect 36070 -5760 36100 -5520
rect 35290 -5850 36100 -5760
rect 35290 -5950 35830 -5850
rect 28700 -6040 35830 -5950
rect 28700 -6280 28780 -6040
rect 29020 -6280 29110 -6040
rect 29350 -6280 29440 -6040
rect 29680 -6280 29770 -6040
rect 30010 -6280 30100 -6040
rect 30340 -6280 30430 -6040
rect 30670 -6280 30760 -6040
rect 31000 -6280 31090 -6040
rect 31330 -6280 31420 -6040
rect 31660 -6280 31750 -6040
rect 31990 -6280 32080 -6040
rect 32320 -6280 32410 -6040
rect 32650 -6280 32740 -6040
rect 32980 -6280 33070 -6040
rect 33310 -6280 33400 -6040
rect 33640 -6280 33730 -6040
rect 33970 -6280 34060 -6040
rect 34300 -6280 34390 -6040
rect 34630 -6280 34720 -6040
rect 34960 -6280 35050 -6040
rect 35290 -6090 35830 -6040
rect 36070 -6090 36100 -5850
rect 35290 -6180 36100 -6090
rect 35290 -6280 35830 -6180
rect 28700 -6420 35830 -6280
rect 36070 -6420 36100 -6180
rect 28700 -6450 36100 -6420
rect 15210 -8570 19530 -8530
rect 15210 -8810 19250 -8570
rect 19490 -8810 19530 -8570
rect 15210 -8850 19530 -8810
rect 15210 -9970 19210 -8850
rect 24480 -9970 27700 -9600
rect 1080 -10340 2680 -10310
rect 1080 -10560 1260 -10340
rect 40 -10580 1260 -10560
rect 1500 -10580 1590 -10340
rect 1830 -10580 1930 -10340
rect 2170 -10580 2260 -10340
rect 2500 -10560 2680 -10340
rect 12220 -10370 13820 -10340
rect 12220 -10560 12400 -10370
rect 2500 -10580 12400 -10560
rect 40 -10610 12400 -10580
rect 12640 -10610 12730 -10370
rect 12970 -10610 13070 -10370
rect 13310 -10610 13400 -10370
rect 13640 -10560 13820 -10370
rect 15210 -10370 27700 -9970
rect 15210 -10560 19210 -10370
rect 13640 -10610 19210 -10560
rect 40 -11360 19210 -10610
rect -6530 -12240 13070 -11680
rect -6530 -12480 2390 -12240
rect 2630 -12480 2720 -12240
rect 2960 -12480 3060 -12240
rect 3300 -12480 3390 -12240
rect 3630 -12480 11270 -12240
rect 11510 -12480 11600 -12240
rect 11840 -12480 11940 -12240
rect 12180 -12480 12270 -12240
rect 12510 -12480 13070 -12240
rect 2210 -12510 3810 -12480
rect 11090 -12510 12690 -12480
rect 15210 -14190 19210 -11360
rect 15210 -14230 19530 -14190
rect 15210 -14470 19250 -14230
rect 19490 -14470 19530 -14230
rect 15210 -14510 19530 -14470
rect 15210 -15860 19210 -14510
rect 24760 -15860 27980 -15460
rect 15210 -16260 27980 -15860
rect 15210 -20260 19210 -16260
rect 15210 -20300 19530 -20260
rect 15210 -20540 19250 -20300
rect 19490 -20540 19530 -20300
rect 15210 -20580 19530 -20540
rect 15210 -21680 19210 -20580
rect 24560 -21680 27780 -21340
rect 15210 -22080 27780 -21680
rect 2210 -22660 3810 -22630
rect 2210 -22670 2390 -22660
rect 1710 -22900 2390 -22670
rect 2630 -22900 2720 -22660
rect 2960 -22900 3060 -22660
rect 3300 -22900 3390 -22660
rect 3630 -22670 3810 -22660
rect 11090 -22660 12690 -22630
rect 11090 -22670 11270 -22660
rect 3630 -22900 11270 -22670
rect 11510 -22900 11600 -22660
rect 11840 -22900 11940 -22660
rect 12180 -22900 12270 -22660
rect 12510 -22670 12690 -22660
rect 15210 -22670 19210 -22080
rect 12510 -22900 19210 -22670
rect 1710 -23470 19210 -22900
use core  core_1
timestamp 1634785440
transform 1 0 7320 0 1 -7060
box -7010 -2490 7580 4060
use core  core_0
timestamp 1634785440
transform 1 0 7320 0 1 2520
box -7010 -2490 7580 4060
use mirror_4  mirror_4_0
timestamp 1634784454
transform 1 0 18540 0 1 -20790
box 850 -570 9240 3290
use mirror_3  mirror_3_0
timestamp 1634770709
transform 1 0 18740 0 1 -14930
box 650 -570 9240 3290
use mirror_1  mirror_1_0
timestamp 1634782873
transform 1 0 18460 0 1 -9070
box 930 -570 9240 3290
use cmfb  cmfb_1
timestamp 1634684585
transform 1 0 23300 0 1 -3610
box -3910 -30 2310 4270
use cmfb  cmfb_0
timestamp 1634684585
transform 1 0 23300 0 1 2690
box -3910 -30 2310 4270
use sf  sf_0
timestamp 1634767319
transform 1 0 12590 0 1 -29850
box -10660 7260 380 17300
<< labels >>
rlabel metal1 13020 40 13020 40 1 s
port 5 n
rlabel metal1 13060 40 13060 40 1 GND
port 7 n
rlabel metal5 17260 7060 17260 7060 1 GND
port 2 n
rlabel metal4 20170 -21100 20170 -21100 1 Vb4_
port 8 n
rlabel metal4 20100 -9380 20100 -9380 1 Vb1_
port 10 n
rlabel metal4 14710 5130 14710 5130 1 Vb2
port 11 n
rlabel metal4 15010 -4700 15010 -4700 1 Vb2
port 11 n
rlabel metal1 19410 4510 19410 4510 1 Vb5
port 14 n
rlabel metal1 19420 -1110 19420 -1110 1 Vb5
port 14 n
rlabel metal5 -2700 7440 -2700 7440 1 VDD
port 1 n
rlabel metal4 7150 21290 7150 21290 1 Iin_p
port 15 n
rlabel metal4 7750 21290 7750 21290 1 Iin_n
port 16 n
rlabel metal3 9730 -23610 9730 -23610 1 Vout_n
port 17 n
rlabel metal3 5150 -23580 5150 -23580 1 Vout_p
port 18 n
rlabel metal4 20620 -15250 20620 -15250 1 Vb3_
port 9 n
rlabel metal4 7700 8030 7700 8030 1 Vinn
rlabel metal4 7160 8030 7160 8030 1 Vinp
rlabel metal3 8330 2730 8330 2730 1 Vop
rlabel metal3 6540 2730 6540 2730 1 Von
rlabel metal2 7400 360 7400 360 1 Vcm1
rlabel metal3 8870 -6850 8870 -6850 1 pre_Vout_n
rlabel metal3 6040 -6890 6040 -6890 1 pre_Vout_p
rlabel metal2 7420 -9350 7420 -9350 1 Vcm2
rlabel metal2 7620 -3520 7620 -3520 1 Vcmfb2
rlabel metal2 7470 6130 7470 6130 1 Vcmfb1
rlabel metal1 19490 4790 19490 4790 1 Vb5
port 14 n
rlabel metal1 19510 -1360 19510 -1360 1 Vb5
port 14 n
rlabel metal5 26700 7420 26700 7420 1 VDD
port 1 n
<< end >>
